PK   �2>Z󁁣d  ��     cirkitFile.json�]oo�6��*���2H���s�{�w�E�k�`wP�5.k���^����v٢<�PN���M��pH�f83I��6�����כp�K��/׫��泏~�|�ϯ���n��ٮo~�����7�ǿ��ow��ן�֫��ި��iQX]�B�&ζM�X���y�fo�5���Q����B�R���`��Fs�l[��ه��{攞�g=��	�ep�H�
ٔ��%EUծ�e�a<�d��;�ٖ!��YQ#�g���kU�o�c�����$�M���-��57����%��_4�d4�yJ���t-(H���I��6jI\0���!-:뉙C�b��S&��i�eZ��6�j^Қ��j�F+�y����mic(X�Ѷ����Ȗ�kO�;'��S�}�t�R]�Vq�m!/)�,l��Y(c��Ò�׵�tM�:'�)O�o��)eF��ղh�iY1VT��Eh������I�Dj;EuM�u��OQ��k�����&��� nk��0"���P��CLdLN���)�j���}SR.1�Ü�{���"6�kR��S��q@��i'�Z��	�	t�P�ZQ�&<&B�)�#16�32;IpoSC&'p���
E)�_S���v�!��g_�U�2F�Iy��X]'�d�=r�?�]=��KK䢲Ȣ�p1Y��,\�nv����e��<�t�U�ԭ��)wҀ�062���A0?al�w��`S��&��6���YÉ��f�rw�Lm.gQ���f�b�Yl&v�8���9���<|y��;?:y:��*�hl�6�m)l�`�����)���A�����Qܶ&��S� �U�"I��"�E3,��a���<(yP,�9C�M����e�E�S(l�l\�����r�}E������������o؄���`�7���.6��hş�#�[����*<l7����sY��Y��,\T.:�������A]&��A/�_��<�y�F�G�\�.7:?B�G���C�G�\����s9�:t~����D�G2�.x������G2�������&�y�<(yP,2��<(yP,�X�A�ȃb��"��Y��#t.g1�Ώй�E0:?B�r�}��G�\·�����5B�G�\��:?r��e����U��,�_��C?/7�����ס�Y�n֛&lfo�֪hk�,��nkVH%��:0UY��u���3'[ëB2�
�U4�⺭M�K�Ǉ�˻攮�]��T�UuѶ���+�^����.�ګ�UHf�oT�<�s�^*^( �)�ua]�0��.���ԘQR�Ɯ�%�$=+�V9_���t��F�B1�/u�J�}�gT�I��je�(k�"LJ�S[]�q�p�tQ��ՊKR�%���5Ř$m	�u�)5e�۝3cU�(/�/*@6��=�-���VU�x]ǜ��gEZ�ԣ�Acuc�Q#� ����hO�oT����(KX�]�i��-���T���V�:�eQV�sr�Q�)�6��s�x�z��;9f
��C:���N(����PH��t]}!�k��*�f����lO�sr��r��IK�<&�R����5e�J�%Q
,&���"�� {M|�k�B��S(���7�Ɓ�3��$ΌwJ�5���H���˶�p�������F�L{���b�Cٵ�����$eCz��Y��6�޶�&�޶�����{NYP��2`��t�����U�5����2�����������A��P=Sv��Jz�����-^ 2ʨ�N{r�2�)�a����=�7��^�A)2 uM�$��9SI�5����Ee[1S���k�9�~ި֔P�6���ؐ�(��TwGqN�	��єw�Pj]>|8T�l§�/���f�*���z�)b�$	�*�I�u���UF�F��dK����x����&�l$3*�5�iF�JM]ji]�eZ�HU6����>�% f�&�l	�dj�-�!�0�CC��G�؞I��V>g��v{��#r��b"Uf��	l�4��1����=gv��T �%��%���% �Nlu�d(�	�
p�S�ivA��gM�5j�K��!L�!`�8'��bN:�5�t���iR�,і8�)"���礮Pi:.�5
��P�N3H@,?����U���Ǳ�v#� 	��w��ۂ�i�瀪��*���Xw:����� �t�. ��wT�k�� �����-@�r�)�s�)L�V6�n�ȑQ��Z_�0x��W�ټZ�b��iK{Gڰq ���8���(t	�1ʨ�U_�Ly�w�)z�-9�"eK>��ӑ% �ّ���tQ�q���!>B�lS�ǉt��r����(�B&� ��:�
�'�h���XC�}�RRLI���>7��C{u�U�)�M|pݾ �D��:|� Ժm�y�T���	��	�P�,;�U�v�P�v&S�3@Q�\���x<�. �)iz�E}XzT��<3�!�$>:�a�OP�W�� �d0�>O��Ǫ3H@|�z�MgH'5�ا�G�����%@!���q{�t�!r���"��ݏJp����)0�C�t���3�i���oi>��>|�4~h�a�P?��z?�T6?eGI�ogܐ�|,��#O�Q&KG�����%�w�әr!�_ݤ��O�KH�j�` �)��)N҄Q�G ���&�ޠ������Oq&F��'����Dx��~_�mRڏ���MJ{���76q���&	�T|r*@9���㿮y����3�G�%�=��m�&ld��c�hD�J"��6��% �W7��Q�VP1.�T3,�vXP���V���T$�����Dԋ��fb|��lf��qM��Û8�G��2Y�6:b?�{��8�ܒ�"a?�y$]�"��9qs��PgFvj@I�����|b�lb���$&晽y7��I\��8�(c4�7#�Z\��[�V��m�B�. �R��7f���Oh��oY��"=�����Ht�c[��B�"��E���>G:��uZh`��)hhL[�ڇBKXNYYUX���B��Y�5��Pb ���`�a�U�F��X�'!A*=��)�4�������!�N��a���8�|��\�����>�&�1�c����4��jR��u�[-a$���B9 ��̠!�����>:A�k�O�L��P��CS���8�ԍ��*ǫO^�6~���W�6:G3}��W��w$���S'���\׬<�'��)�ý�[zK���[���A�S9��v���-��eOo��-w:0~?mv��.t�7�&��Z�M|�z���]�ow~_���2���oc�{w��f}6�e��Ow��_��y��,W?�<+�)���g��ۇ�ן����Շ�:��o�ן�[}|goZ{��}����_V����&��a�	���v�`P������a���9�3I���u��f�D�[�/��5�ûB0�pJ+���T�y�� Et	s��x�Lj��)����R�:�o6��,C����_ջ6��o>[o��x~'��6�q��rS߆���+�1��X�3�c����0:�RK#���0�-0@��sh�0V0�����t��Z��%�t�\Δb�K��Ǖ\8-�0;Y��s3���6C����Ʀ�X��n��Y��O�~F'W#������q� Xuh=�B��sc�C��t2���'3<�9��f߫8��F>��:��3z?^#���N:��df��������t���=3=Lv:�b�����}h����~g��hݨ6�t�����4��<,�_}�jbH~��Z)�-�Ԃ��� �疩jJ���N�s`�F��	��k���h�Uǖ	�:�L���L���o�伴,G8�`�K��7^����`��,w�A΅�Is���ϐ�%��q�'	�v銪Sn��ං.�*v<Cw'�#��(0Ij�w@`~dYv����}01�	�����+�^����{Y�,� +�����.L�9+-� Y	���f/Uit�v�w�d��|4lXrwM%fKظ��R�3t:n1B��֞"�0iL���.1\!`�`��Y2����`��&�fO(�%�u�sm�~����Js�b���J%�oGŵT��;���Į>L�S��� xR`�����c�� ���sئ3L�)�e�T#T3�8yP� Ʋf{� ��R�Q*m7��{,�� -���Q��g>�Lx��>��To�)�=8LsЋhOK+��ц�ҵ�,Jߺ��:���,D��(̫��QTv����,|_[t7Oba�(���\j� L�����q�y��q�7��+t�.�����D�N���� �ۣ7ɘ�����c"��j/�r|� Q{�ϗ4A��%�u!k���-�g��y�Gu6r�|����t#,��)�])�b~���,�SϖvG�"�\�O ш�w�xr��~��_����}����yu'N����o��ߞ������+�b�>�+�;������7�����i������HS���?o�������W�$�1�Ө�n���?5������ur�z속������Ow�I�Cȸ��z��a��0����#S1.dl���L�o�����>��wd���������98�`#G��J��~p
������hx%lYh�z�^e{�˨���.m�]/�a�q5�@:;0�Cl�s�a�j�a�Q�7<>ykkS�qWW]��'���P<��J�) �1qC�87m1�U�3_�5���5_�\d�'µR)حM��y�l?�[�p�9�kC7�x)�c��㖿����_͟��o7a����e��S��cLJ��V�������ת����g��`[����ۦ����YX5���'�����CNـ�_2�w�^�]�ۏ��߿?�i��ڷ��ݎu��y��J7��!̇�y$ףz��a�_�Ͼ R��޶�}�#O���/�%��Zu��E?^����[Nv��{�,U��~�zʀ�K��T94��Z��@C�WߑgX�] ݥ0{<9����҇��OQ� YL
>AMf��V�jۼV�����e�0�-E}��nP����2,8��~F���|[���p�u��/�G?���K�����Qb�*â_0��W���"����.��i�r��$PT'[Ej�a(&�����G�Y�]V-ߋw��O`Rj~Du8�}��wWO�2(9�����
L��_ b�/�b�~H�w��Or?��}*>��3�T��?4p�������0��7���'������'G���h3lfd��6þ�C���t�Շ��-'�j�f�OS�TX��Z �ջ�~.�n"����p@*M/���:�,{�秓�؟K�2����My��/sS����5p�1+�'4PTO%����	U ]0�Y"�܉���#F�Ë�[�#��$hw�8B4��tۆ��ȧ�2�Kh\\"ޥv�W�ry����X�����K��"�˛;Y�!^d3���F�qD5���)�Txh0Ys�:�7���~/[.w�Eg�O����PI'C������:�Vy���$c�sA
��rA�E9�~�w}�Tt+*/_�`U��^�!�|�en{ Љ�Ļ���W�Z�c�ḣ��G��/c�������o~6K{?{�r����wh��W��O�O�nç�8�_f_�PK   �S;Z�%�W�  ��  /   images/538bc4a9-05ab-4361-a8c5-43654019cbf3.jpg�eT\��.�$8����;��{p��=	�ݵ	��4��ָ���s������8���=���=k��i��֜UO��ٗ�8 �� "" "� !�~����-2
&:&:&�;"<lL<r|bbRRR,����$�D$�$�X�5	6&6��� 2�ޟ��
�@� �����W���������O��/� Tx8�+Lx�?+���p�H_ ������YH � ���?� �[y���g���N�[)���J�!�j���m��z�۝�iJ_ޫ�^o��mg	/ʽ`q��r����'� ���G{�U2�p�tDR�`Z���f���������~�z~��������Zn�ԛ��7�E�$	]+���pr�6�w��`���%�Y��tu�	,�T�$H(���.��*����wIb�0����@I���L��f�/M�k�e^t�;�כ�'QS	ʳ��
��:C*�7g�C��e3E�4�@��x��Ψ��������k2 ��LH#��H�bf��,J���b���G��h�j�g�m�WD������c����<:�k�:�x07��b/���I2�;��U��*|��?"��<=��$A�s��H��'�����#Ir}�·�^�ԟ����7np��&S(Ҕ�7���~ߚ��v��I����vy�iCO�vY=*]굾��"�����-��%��p�{Е�i7z��]�'��ϔ�jk2$��̹�lk�����6Mh?P_��2~͖��ZDw���Y'�Â��{¿Fɛ�H�lD������t�ϼ%'R#g� ���t�����}���N��J�]]��=u?���P��O�(�u���YV�{Cdt�g��
�X|�|�X����R�C3x(VI��(����ZF�X#�SI�s��Z���,�L_�ȉ6���G�+�9��"����Z�f\^ri�ܾr�m��`�>����WX_��"s����7h#�
�-�]����ؓy<6�V�:[��m��"|m+�sD ��hI%��_3A��s?�z�!a��FE�
���yxn�N��蛭d��� �w3}KW��(��4����0���;��g�ϒ2�R�6�C�cM?�+�=������U���A�@����4�Q	ׅ��l�е�,�?��ٳ@��ȥ�˟	���)��Jn���
ȿʹ���4u,�ÍI���9�벵C6��h�e}Ym�X�w�OF��Roެx�7��7��D�7�)>hqy��>��Kq)�y�n��FZ��԰dl���n��[���b����\e�v����p"�	҈a)c^*��B�'�  l|"`M6J�@�WA�vs��r��jҒ�Yԗ���-����.��(d�h�xb���He����2��<�������;*����q��ff��'��Ɍ�j���M�o��l�Xh��0�������Y���J��:ؗ�2�n��:Q�>euf���#�%��S�#Yy�����M5�fp�G���4a&�kk/�K9uf>�,.R���v5�Z�^�����K0�i^Fցmm8�˪Љ�3p��Af% 9uP��y�.NM�)䫝����z/�}�F�t"bj4dg�I�i�e�׷rJ'�b[HtH_$����SCV�M7����_Ӭ�XB��mB�2�E��n2@F�Q+IvO�Y�7�#���f��
���{��"�c�7,�X]�xN"��k���«���w�7!�ʓ����ΫTa�����t;�1|���e�S�Ӥ{iU}��%E,�D&���.QN��A� �����"�B�
�ſ(����7�4K�5M�X�\~U�fI�r�-��U `�S�$�E��c���l%G���8�����5�40�U�����[Ɩ�I�ਔI霺��Q��NgmO�ʥ���e����MWV��r�1 ~��ۍJ�5?[Z�)��ቿ�ZXW�<��[�Q�,����s��Ʌ����e��_����36���%|��>��;t��:��M�t�ઙ���y�ƠS������XK�D��Rq��G��I��c��~�[\�<�1Ԥ-�v���)�ƃ�MU3�	$
U�`͚\r��'�V�o��ڽ-|���J<�̕�M&�0F<�K�5��2�\�_o�>{W��9��]�ֶ����d.����e�N��Vx�2��ra	o��3���$��]L���>��6�p��z���Sط^�ъO�0����湡 �_,K���9�[�"z=�Ku8U���L�[���Ks�㰋��ǻe���~Ϻ����ց��c/C�e����A�L5�.{����C�!����Ҹ~e1� ]
���Dѝ�����Q��{�t~$�fA��}�u-�&韔 ��
��tP�lT�����B���B oj>}}�n��p�x�p�����S$4x��&ߣ$��]�f�ѣ�f(��!�p��=0d�f+��aa�i㡄����$t�0{�)���XO^|ѪۖJ#����g�5�K�(f�c&oT����P�2~���v؎c+^Y��p�Q�OBV#;a�ۘ���j4y�NW5�Yre�Y�\dv��//���9s���_��fm'����o@{Z�m}~���Z�-��$��r��^Y~袟��|/F�I~!Ɣ���)�^�ܟb��"r�����RW-�ibN���1�� |�Q�,��DF1�RM��s�C����|RA��>�q�=Wq}�7�HE� �3R�������[�^���G4&]-����~��޲��*��9�rq�NؠYW�K�KA�T��pb�!�`���%���J��}b����3��Ǐ	^�@�W�$���C7w�ۆ^�H��Q)�K[��>����Ǌw���	 	�7���4J��GH�S���b�h���o���9�룲S_ �Dʵ�מUG�XX��/��؃�'���?�=3�П���F�Bz����[�@S�ד�i6��M�f9����~�2?����y�[z�O����PgȽ���7?��,�Bn��n�|Yǭu���Hak���dF?�r�(�;�p�j8N3/n���m q�<L�hG�����8����<�B0ѱ,��߉�� %ZYZ{l��~�.L,U0R�����4|޳�}}�J��L7��_.wA*�E�Z�oֵk���cՊ4!��9���=��-�R�n�^�<z�U����p���Jt^;t�{B���.���K��dS>�,	۳ȟ�8�qd�0�8��\�g�O�6S��s�PԦ�3�����v`FB��i�`���N�9�_�d�wW��I,�*o�Rc����Q�k��c�`��4�'��!$+�6EW�6�����8����������Ɂ@$��⍕}g���a@&*�	&�F_$��bՓk���l�g�4f�S��r�`9�w4ƾ��w|���4��Y�2�D���%�|u�`�r饱_(W�&�K�i���+˘5O>������f
ʝ˚�6�����i�T!�bi�''��ǻS�nP4��ȀϞ�v'C(F
�����K䃭��?��Z�Z�F!ֱ��!v[���l�m�p���U�|I�"��#t�t�P]O��|{Q�gڊ#v��x��u�陵�2��T��:vX�Â4�{XU�%A׵�,��U��������+��8p	^�|��{�c�h�FU{T"�\^/n�o�i�PmPZ�ۉ0\ZomY�˄��s�m)&x>d3z>�7.�ݡ�a� >:��CM�M�<V����,*#�]��X�뎙���_6��K<�wdV�Z�':�K2dd�DiK?n�f8�\	j_%nw�
XǗ�=> �٘�B��J�<x�t����J�fnd�1zB���6��r?x�K�'���)�%[��Jk�y=u�r����9�z�7������~�KG���dw�gp��V��3r�y*2~dɖЙ���.Ũ۳)�P��n�	��[>H�ގ=���C���4�G�K��M���A<$T��-�5m���ܤe"�-���Šq��{9s�8����|j�'���Z���A�by�q��a`M��� ��t���B���g<L��,j�[��_0gN$�$[L���4���(Ѯ3�'v����6q���5�魞�|A�`���4�w���p�D�ĸ�e��$��u�����t��6�
Bid1+iZ��Ql�W��h�!��ut>�����C�Y�ͭ2�[����o��`f:�ዐ�G��O��ޗ�O�����c9'����h.�m��W���(מ�6��4�$�8�����=.��[� ܁J!!!�)~u+HA(�qPj�j�bU-��ɝ9so�g���^x�����g�u;�!;_e6��C��Ap(٩���7QBac391�K2?�]G@W�'�q�u
�&m�^��7}u+y9���9����R���;Ԃ�Ps�l~��ֱ&.[!��2}��e��Bv/)Hق�������6��RfHK�屒pη�dk��J����a�:�������=mlQ�p�\R�ƈ�Hs-䠧<�e��2���@;'�Z,��{,�W8d���vgڂ�U��'$iF���65Q<Z8YǓ���,jHg��;�Wb\�Ed(y�jd�r\ג6��_M��6��<v�����%�;W��s��=p�c��Yz:;A��{�5*��Q����Tɾ���k�A�T����m�~}����a�{�r���.���`@ ���!G��9��j� 4���`�t'og�S:>������eQ��!��b�F�+��W�Ņ٣�v�m�t����ױ���=c����"�~�v�{k��)ޘ�&$^�T�P_&:�@��2� �rb�Ǫ�MH�%�%Lo���k�Wszk/��b�=C��E�?�װ�kV ������\�]���9�!:/���)D�b���'e���@����.CM��E�����N�e���H� �#S��[WUqo��d j�Z�h��	u���r����f��f�\��ψ�%���4��zx��B��pYܒ�{$�a��m�;w�߹���[9� 5TVS�f��[l�����+�y�	�W���m.�˪�N����:d<`k�.�#�����P��o>*y����4�Y�~�8��>�J~sb�X���-!m%��^)v����z�pa>o�.s��X�8����@�rM�����0V��_&�'Fk����'<�8�|��r\2Qw��f��T��vlwj�]���|��I��C�9�M�WH�[5H�N�|�2�lR���%������F��Q~��CɫJ���F3�FJ��^�آ��+:mj�DHn�� \0���2����?O��N�l�n��[|�0[��~��&���!_�� ��8G���
�ǧm|1��勩:Ϳ>;�.!��R��S!��!c�!�#S�¢4�4�����㱕}5`�b����E�㣤S��4�_�b=@N6�@�M^j�+�!�&�0z�����Y1FA�̙����'�$3�
M9��X	��� ~��\XfjP|�W�.#�V�!l��C�&���'b���e����|S�ܸ�
1���w�J�B��(�b'zXc�婍�,�.z8��9��K�	<�&�M2ξ���?mߒD{
l�H^F̴�gs���R�
 �#T!K�8����{��N� �;�5��xC��\cu�覰,-Ԧ�Ҵ��r�9#�K�{����ɭ!n���t�a���'��0�"���$��/�sy�F��B�f!Y�1��8ZQb����A�i]G��H�.�O���9B3���9��Ɵ�CG��G�q��4��1���~3������}ZH��O%c�{5�^k<h�ɉ ���)��m�t+w�ï�<�&g��)bs�-��-$Ԏ6WX�!���	A�NǺ=��j��O�3/)�%���6���-�B(|�Z��C��I���o6Q�߶�_R�eL">a� P�r))�֥�ŰB��҅(�"�$���E�c�y�M�Օ��f�T3��N�.x����s�������vv�����r4���8G x��W�E�ٌ�C�!+����&��(�W���_��(hD��!�q*��m��>`N+Q���f�~[����T��?E�^Q�+U��������:Χ�s��a2BS4�d�� Q�b�Ob8�To�)�%��w��A���0���C1�ƪ{����BQ��'�׍��k�*�7j�x�0?3L$�1g�����Ǥ�)e�������[6��(��ϢX�
���cR���F�I �꣢a���W��ޙ�O�#���hY��M�,�����i�r��i둩r���#->�ߓ|��]Kop ,��m��#�����©[�[Dg֐����|�a�S�P��Y9���B�Y�i�۞�E-���#�f��
Yx�%�'�O�1�~gA�`J��k�8U\�G�`�r�c�(i����u��:w��F=^�[�C_�Dڸ�4�����.�8wM���`3�!��ۿu+o7~+n�(ޖ��,��vgŗ`��9ށ)��P��Qlӓ7AQr1I�9��{\[��\	��\��e�R�hJ�2Z6h�D��-��cu=�E5����p�f��rR�h<���R���!���D�vm
BK��͜Sh�\ЀT���o��vҴ����,i��LS)]����_�k�����_�o�������࿵��[����V/] NL <�kDx���7
8�+x��X�8��p�(>��dcW�������d$V)�2@�3����m�/�@O����������Ђu�r�;������O1�Ks��m]Ѣ�$�|�����[T�(�N5�0�PWy����%dȺ��{ھ�� �^{{d���������r��7�5�	�HD�"P'���� lMe�O_w[A�e���Q� 3��<S�q��m�'9���=-c��9�:�Gy���6�([@A��y�ps���%���I�B⡈���k�#���[�Yvq@l٪�g�Y�� �'�þP�U6
��O̧��bGm[9�~� \ORqAq:���R�Z�Ƅ�����o���\'ɼ�3����Y)� .j�^3��v#�z�
]2Y���j
}����3�D���OY�n0[����>�m��"��0icőQt Yb-+U4|��{�W �oИ2�w!A�,�������#��#��uC����/Sm��'���������(�E�ٷҜ`>���9P�l�����p�ձ)�֗��V�����$w��_R��LA{P�7��uЍ�3��^(��|�ލnln�`JaS<�Ք��*r|�$�������&��6���ft�ML*���ش}�>a$�i�>�[ߤ�o:pb���؂8�R�4��R��V�E6ހ�؄ب�,�����è��p�Ƣ��!4yy,f�9�_��'I.�K�|��pd�mi1����g��f��Ս���8V��`�V�w��}�ZW'ժ��	?����UC�I�����L�K�䒓�M�@�����s�з�V�LS緈���oV[����|y]֝Urf�%nH�
�P�`]
�o oO��#U�0�P��( �\���$l�P	w�͊�٢�U�^��J���Չˌ�W�|hr����s��͸��a �viD�w&�f�9�&�Av��,�i��W溏X5)�{;��g* �y��L�w���J(��L�҃�h�.,��V>^w,!E���ƐB��//��<Y%v�Q�Q�f��;���wB�?�Z=�rb�?���CW]{lPS��?-s��g�c����uJ�v�<�?�	&��NS���Z	�N��B�1�r�(�����+�D�O���\ڍQy$�3�-vH���S�b�Wd;��l��Li��ޟ
�2��/6hB�;��w
�j2��/�?g��̓�}>��q{7�'�zr���J��r��tg�uĹ(�%4~��[8��Bj\]�w��VB�l���?�2��S@s.��jS	߮lv�DwS�82",e�
&���Y��(�B���}�r�S������"4���u����ů��Y�B�����N��?�q�((��n�Û^���/ ��xOCv�$s�����4�1H p� _k���| Vx�����1LǒC�a�X�LĐ��!�b� ���#>��^��H������5ޑ�b�;��V�S�2��:��&ҭ['��ɰ�Ǉn@�`�Ǣd����&ir}����]P.^���A����&����� A��� �6�E���V̈��}'����p�i��Ttd�@� ��AM��h0��ITi�E�=�z�U��~_���D�k��T:���Kʊ)i��˵��hj�pB lz�^ŧ�up|sg�Bj�c��?W y��{���x�xB���Z��k�B�nI�h��h��ҴO���R��a��� .8�?�i��xu�7��������R%�k��Wn,��rJ�W���,v)��T�<��T+ħ������=L�����<o��l�x S�@%����� �o�=~�0LU-t�ZC<+��$�^��ԌW�K��WR5	jQf�V���v��S�v"�$��Z�9��qJs#�z-V�b�s ���c̉�>U	u��A%�J��t�*Қp�ܯ���_��)���P���p�t^�aO_>O�y�ԡI��`j��Ћ���r��&��Yb�5�ғ[<��4�׀�+���7�W[�}�D�B9^��&>�>���k�f��_�&�sH���O����J:�����_f��59�ꅷ���b�@J�sG�����n��5��L��X��*�K����Sw����7�8br���v�l^����	���l��\��X	���;֑�c��.*h6-���^�bUe�e���b��� �.��������H��F��}Y�Օ�[g��+l�,�~���*��Bl��]�OO~�������3*���XD�ThP�����Z��n�e)�w���3�%�<Q	����=Z��h:L4�ng��-�:H7?.��:��o9��aL��ߓgݯ��M�r�/~��15ܢg�p�ʝ�:xk�N�d�.|���n8���B�\��(]m�xe-����j�T�<�>D&T0nq���8+�2maM�i���C"��)4}V@�JL�^��e^�z�b$ �g�y� �7�/������a�t��S��am�xo�����\ם�b�(�����#��Z@R ��Δ��Qoz @���c�9%����"'zX��N\�K�5���q�:�Q�-�r�Em谾t��a#�P�h�w�|q��RfE��F��z��T4��
�-����dU�ո��lk���p�v���(�a#�sכ� ���!�}4�Ih�͍����{�ma�^'����.��ie��%��ֿ@פg̑d��O�[�M�H^s���aK7��Φn���y@����	a��&3���˴�]�4w��ė ��v!1�?�uǬ]6hI~�"{����u�'�3TA�jBy��}��'�	�
����N?��<���ӟ\v�9�}��9�L������1Y���r>.�շ�g�aB�F�I`�f;z��d�wacF}�>AΝu���<�To`�$EoJ��`��������$�i��ZG�K� !�����Փ��r�N� ]�zF����1ټ *�u�P��0���92��IWA4��%xDx�p�}�����Z��Ԍ�E���N7�[ꤤ�f�"�P:�^���7�����X{R�����?-n�j�s���_�����͎5�O������H$�qKP-��y�p@��߭�q0v���&�Fd���-���Z	O	��~8
t
�E4?g�y�1�y'��PlL���!����g׬�	�gU�V<���_����>nU|Pȣ��:����!f2���8o/ǾP7�P�bS�=e�=��ܻf���KJ�F���/!S���i��]�Dm�klUm��������0^���;�q��(г��0�h�<��:�e�X͎�{7
���@�c��V�)���Vv��'/R�44��?���X�*�ȉ�+Xք@x�ӾmA� �X�2����G
\=��;����qPh>���=�Ȧ��4E(�Ý�K��?�<�������NE�
�Aj��eD�G���7��#�'��J��H�%��}F���E�pXd��ϸ7	��Z�`�8s*��y8�"P�Z�+QC���\���`h���w��)�8~Xdtk����{��3�0�)K�*u���;���v>i>��9o�dx"��qˣ��5��}6_^��D�����MT!Myf�F/�k.�+�,��)�ſ	�� �㎠�ѷ�=���H�ι�T�!�K�9����?���ǖ������Ҽ�W�F�5�EktE���a���.īU1#K�_td����M���]��킕���vE&u잼^�s�5�E1Z���Cy�>@~H����Z�VDe�ј0��$�K�u��wo�c���QeSȤH��2Z�<X���6��S0##�*�6����n�Jɘk%��)��g-�%���<��R���F�M��7�C�
��*]),~�׋vK?��u_�K���Ť8��f�_��x�p4��u�Q1�K�G��U�l���j7� �i��fPM�ͷ�����L��ڋ�Du��e1Re|�XB���{�-D�X�s�2'���B���`�uWe�9��u�ӟ���Ƽ���������)V�q���Ox��k��ӊ��Q@����� /�����/~P���%1~Au��jWv��T���/��6~����6hK]��b�v�_N�Hz»���Sb�=k���1z��Z�M�E���_��r��#��h+-O��(�G��F�:4���N��	I~7�������������������l�(�#���ȹ7�cP�z?IA��~��m�KQ�'|����3�0.`�w���/������&0Ŗ�A�ڷ��Y�a���,Qxh����P��x�[�|2ᦛѕ����p���g_������$���hr�e*IdQ4=��X�\XK^J{t�;�Vo�����;��Ď����M��^����ih{Ê�uL�Qo�ب/��d��\��@��v�.ƍ�?�(^um)�&~��?�66Y�`��8	�We Gdx���MF��C:j4*��5$4����YK��v)��x+$��Bɯ7$g}>�Vn��HoK�Tf��g9Y�Ŕ��<@�rR��.b���(y��)����)�`�k+Ao
�U4�i-�����\��������B������z�o梏���;]j	)�L�M�FW��U�_��ȿK��MX�뢫��O̓V{r�h��-s���J���g���~:������u�X����e���}��2I��Q��<�%~G����O���W�;p!w��K�C:�MC=��7F��,~5�~�`T�yP}d�^=�;�RB|z�<%"
�(/֨����n���Z������z�Y�Dp�b��|���DUEn� �I<��zؑ�S���Q��V�*��r�m��K�gD<d?�CzZG�D�	Cc�M ]�x�U:]��DA��/ {���}�g��|)OCjx|������&/]��f�k��Ԯ�����㍼ࢨCI�0�ќ���l�Qz ��m3���"�xuk2e�<9�W�������Q�B��5�;�ڊ���l�)����o��:��c���;�u�l�����ȏr״��f�g-���Jn�+��ww���9�֧Ր[�[eP�:�e��`��ۀ���AO��z;�1��n�����mo�T�/�)��G}h+�T�&��Z=�vq�PԜ&�iu�0�>����T>D���J* "ʂ=�`\u�FB�����aL�	�������fƸA1��'L`f/E�f��=e�k��g�#�d�CD�̹d��Qr̕��'�9{`~�V�+������������`�>+na�d��s��1���F0/���O>[���aHToJ�L�A��g�v�\�ǌ��_�؆�!��ku��;�e-
g�X��L�>'��2��es��wx$!g�����>�(���F>�Q��_�DL6,+�OX�݌�ݤ����y�Jڹ��7��脻}�#_�ĥ �MLήW᧩qI�4L��J���*�*q�<��b󇯩�AF}�!g[Y`���gFE���#���mN���9{$Uig=!�Dn=�ɨ3������AR��Sl��gȷJ�����/}��;@h7�1������^�ʿ�>��Tu�M�f���eݰ>Y>�^�Pz,^K�h\���h/B�����oO�s�k'T�:Ϧsc�D��̚:~���X��}I'��_�.�ٴz�S����^r��1�,=��b춍� V�ݯ��^�LX1���ݾD=�<�Aj�Ĵ��;\T��^:1�:� i3F�荶Sr�Չ��z1,T<������%(��|ܾXΦ�}q��U[�"`��;:7rg�:p�dB!�刦tǾ ^&�}�DB�cL��E���j�٠� ����}X*1��oM����������&����vw�䝓��iqɟ�du
���/�
��HH�V�n�V(����x|�y������xV:��������w�@h�B�ԭ���vo�`�%�g����	V}��[���I�R���L�5nߛߏrpR���"0�;�s�Y��A�w2SB����.�}���1g�0є4�Bl�~:��_v�#Mt�8I_�	�#��_��q�Uzi�e	/�O��/��~z0/�s(\�.��N�}~�����6�] �ã�}��
���]jbN���t6�w �>�MS
']f(����M�z�fIU�k�v0S�6��,~�\�5G�[�0}u���R���o8��]�2�5�rSp�![Jz���߲ǻ�1�N������v���P0������ V2���/45I vh��pV^cH4wX�Ǳ�m�kF�݉�eO���[�L�ؓ� �^��K}W�7y3c�!�hG��O ����$��Yj��[�Cƶu��g{�De��HA��!�Ȅ�����"�J�����J��{��� uS�f��z;���AJ]�V��Ó>���p���-��D��n��u�3/ �f�s��K������3������܈�Fs��^��~ȟmiF5�#hw��e?��=V���ϧ����~0�;3Xd����O/������8�q!�ր�����La4���Ͳ
����4��D�,ѷU���V>)v%E!��� az��F�<��N��Q���b�擳�Ҋ�@$�����ي����/ߧV�c\��L\l�	J V��д(�,�)�l�{;����X6�j��\?�J�Ȋ=�./ԨVkV���%4�n-����{ť��Qٍu/O�5�K��v���%n�Z�-[��q.����\��^��eIٗ��/�:�1��ɹn�4V'�[�Ootr^ �S��?^ ��G�������g�/����}+��]�)�$ejQ��+�@U��Ɉ��&�v�Șp�D��$jI5���I��jb���R�gg%4Cp�����^��^���h$�Mjs�F�j���]2�>�d9��^`s��%ޭm�Oܟ���J{�0�z���x�j�}7;S+C�!Lj�ǘ8��6���~.�OxQ_��� s�y�ы�W/[H&]�o(O�mlTC�b��ĥ,��Kr�Y+�W[S��k�6� ���fj��VN��^�Ȣ�p�+ Xz��ۏg,��o�|�����Nb���,�eA��g��]$�,�.-��N��D��r�d�$�mV�9��$�$y��]ߪ�$�V����_u�ͷrk�
g�Gf�$��g�T�G�C�9ݗi����,�(���ӝ��SV���8�gWSW����H�ǥ����OЫ߹��8^|&��A���,�� +�߈,C���.�^9������<䚴���8?��u^C�;\9[�'��o]��RRJ�B�i:�S�+|�7�$��E��hg{�I�n��	^<�O�<��B�H�gKPL碚�;pZ<5�ې��,7X��g�+{xmdЭ���l���Y�^ �n�:�EI�l8��cc{sZ��6�TlsG��tVZLj�`���.G�g��z�x�j��
Ǐ[څZ�U~n搙�P��I_�B�������N�ᴒ���7�͔i�6�\
�K2�L	V��M_ UW��Rgh2��7�{_:�Fa�rKg`]��nfG#F��l�[��N��qo�|��:L�j[�:n✫X�����c/��U��r�mOk|� 씳��=ay�8ߣ�$_?Da��?��`47>���:$��֩���2*�K0;:��K��6cR!��I*�)�	�	��)H���QH~�6=����9��E��R׳�)�3A?(�B)��S���y���^�%����w6��/���.�a��=VE�� �YWJs������������a�˹S?}�}X�"׫�{���$�5���A�o�qߝ�&a��W���0�xvWvX�1�3B�M3T*egZ���٥Ae�Ɓ�E��SϼK��\��<���H-����p���-���?���*��uf7��6��Tx6���l�W6�fx�W��j񑐒-skc{U��[�CS&��S�(��-+�z
�g;���qX�{���Ҥ8����^c�9����[~n�l~�<&V�
�&1�-��
��F=~"KӲ�NKK����|[����)�@����?	�'h�0���Lu��{��I?t�K!>�X���
�ګ��HN�e�%D/T<����Y�k`_�%�֯���*��3n�D��&�8���.��`|�%ZQ:f&剤�@���t�H��۬+�1F��ފ֚�Z�טV����dFf����N�@���A���O	B߼T.���\W�,�Ȥjq�-vj����|}J��De6,X�ѡ8�-\'U�=p�o��~P�+>�<��rA����|����h	�5l+�t�������1�6���"�[#H�(V�k�Az�i%*�J���4�yD�"X��%�M}�&IqPQ��\<9�*se�#ŸO&�^�G������5�v֮�6tj<���E_E~��:���۠�]�q!�=�m��8��_pB�,i�v����ⱐ$?��$X8�mX/^Vs��zk�w=�����V�ig�8�F�S�»��}|@�}L�_)	eV��:>��=����0f@K�m��s"��{$�Y0�g�v����,���s"��3cj�`�Q��Q�5����0�F�����\ �*0pC���A���.�QF���M%��TJs��]�E�F��.�f묔�ilA�%�K9ޕNc����W.7i�b��FeX��҅��Իi�����J)��n�Sٳ
#a�2���9��DJR�o !/S�:��_`N������p�M:�Bl�	W��V�\��*rh���:ׂ�r-���4����>w�����'f�`��xg�놽g��u��2��aM/[�J��a�^ʓ��8��;��L��Zl�[X�� C���]=&�Gl����dJmK��#��Q���k&I�$$��A�rh�﵀���n�@�j��RH�p�����9%y*nG�wi>CC�ђlf_��<�g$k�q��@���e�>G�J��sFX
�\	�G��U���n�m:����^�k�Ӈm��)�0������ƅ�˹���b�pM62�vTBkr�c���{���$�q������I��c?-�-���d�V��:�w�N.^���}�d��������Nn�?N���	m���n�������|Y�&g %w»*={�Υ.D�WpC��T�&�[�+��K��DJ�r��%6C�m�/�6��k����]	�x��Qf��f��TՎ:��vJH=���p��A_=sf��A�#̰]߷�ȊL"�5gM��<�d� yYK�e�Q�2c�=+��Z�wx���Xx��E�Y�Y��~���y`����+�~�}���M���Qr�oM�N�@(�#�� �]MR'nJ"��!?P7qECd���y|�XNq���y m�3�E#������~-'��zJ)�e�S)a9^�K���[W����M���~��v���k:��,.eu�?��	��^ ���716�|8wN�y��}^ �_�n���\�<�w�,�g�\��Im�Q0��2{��.Dj�����+u����:[3��4ڶ�#�%��|�&n��u��(D���'M�o�8�{��$�Y?`8���Q<�;ش��6���R�l��MH�ɱ�>M��3�`��ݞ��Y�Ȱ�g<�$,<�i=fzX��)%�[�+Q�:/KST�z�Q�}�ce^vt���X� ơ�����iO���,Q�O;�ς�/*���>�9�j��a�O�5c�[��ǀﳣ�_�˿���r�![��/
^u6��x-ܝ��Bql@����̾4Ȁz���.�͉j��"m�u��z//o���!����b���ϔ�p��+
�@CKs=�,�͵���>�1�P���_�a�_���g�pf��*��|��q�R�2�`~�r�^r��R�f�+�G��*�(�&����=0��[p���������&�w��.IH���}���U�t����u��ޫj����*O<:l��u�`Y2���t�	;d��f5;L�6�U5+~k�W�M�aK�'v �붎,ِ�Հ�.�G��3�z�`��B���UP'j��3<-V�wzs�
��	3X����Y�'�xnE��~��N�B8N��_�GgKc��e�lW��"No1e���s�|yx���5���}��������7lϺ���!�O^��S��[�N�#���D�?W��ru�`��v���R9᯸�����M�aFrp�)�;r�FvS�l���θ�î������"'�1$�0ӓЂ�}�.��e+�E3���'�Z�EH��Rh�w��{�ݣU����N�\e��N߱'��U��5h2|��(Y���2=tR>c}�-c�L!6#[í��s�KG�k���4[�	������g���JFȫ>q>�:^Q>�	=z�^[{FX9h�����a =6  ���*8�`c�R�P�s���J�å��O��b0� �3+����un�_6����>]��)��Y�xHH}���Oؒ�{�W��L�+[�P=�U��z�3�Ɗ0Ǌ��S$�8 {�V�hI�0��5�Y�:-]���HMr��;s�Z�����?�����[;W�G��H�&�L�1�n|_z��a���|W�U�bp�c泶� 8�;�.��禍�h�4���r6eM�{FE^I�>�5O��n �x �X�z�F��
ß����h���*�Pm��
F���3֞Ӻ��Q���`�Β��3zP�����qҮ@k�/}������tn�YW���I���}%07K`��aZ��B��*�z̫�ݰ7�D�$�-�ײ��f����1��Pfs��`�J�-�$ߘ��S�v��W:�X�M�/�˧Q�4Ы(-c�5��B�vv�v���aP�g�:l��kDףSy��{2iزL���+�]���l\y�ᒫ=?:Ϣ�uu�������vɹP�.HP�(o'����K���ȿ�v�@���HW�ųm�'���h�Bܵy����	�ÝHV���H1ߞ}��_��f��l��)�������Ft'YN�n�i�X14iȱ�/$��	 �􏆰p���@X,8��((����+��Q�?
���*�V5�i∍f�~ER4�Q���o���ҵ��}������2+��ˮ�eǬ����jG�onU,h�Ps����*�T�ۆ���3!�6W9�z�B��ztjѣ����1��1o�p����� ��J�J^y�y�t�O� =����������?�F�VL�1l�\�F�Xd��j����X����5�=�I�DKc8�NuS|q��h����*d8����ؙ��y��@®�jP5O˃����N+$��r�� �{�.S�jP�����(���J~������B`�B�S}s{	'կ�4N�g^lɨ!Ͱ��/��,�X/��yRu_�J|/O�`u�c�ѷܨ��$i�iV%	=�Rԯy������!�����l�T:f;%�X�p��,�ឪv�\���Ͻm �95�MP��oa��(,
�a~�j%H��,<�6s��T+<�و�)�c��\3?�j��
g��1rb+��A8TgC5Ү+�u�/���|���p��ƚ�����4�>J�mϖ��57���=d=ٔUJX��@�2 g#�y���=,���6��(A��Ǣ�]V���m���E���)�����P.W�U��]��h^����sG-
>����������u-����+����m�����c���&��3�89�	xw}n�x��;��z_����o��U��;&%=�lB�L����ȍ�﯏w^�)�~ٽ�y?��l�_���FN,��@���J���8O�6)aKK�35��R���س�C�I�GB@�������Drlx*,\jN.	uJv3�4nqI5�0<s�ZS)��f|����M)G�}�]�h�wK�@���F�lY*��db^s�i~�< M�3�O���Lp2|Zп���weS�S���@�O�gY���e .Oq"�CY��X:�_��o���1��MG|Zr՞��>h�s�bq�{��L���$f��ɜ�ҿ��{��u��d�Q��\y�&'�$K@��y�3VM�jSn	��v��"�/r��c�f�c^�UD�IS��k�WVؾ3�a��G��&xL-��j	x͇���L^�pV�u�/3W���W(��I�En�]�]P;��Yam�,h�rк�fp�Xv��'�b&�����խ܏\�R\�8���O)c���6Y�w�*�|d�t�_h����7���wʱ�̋3}d��s���c�����(&���w����`�<w�O�K��N��y��[��y���uw?Sbm�XԈ�`I�i3��}0ʳ��,���G�V�y?�!:� � 	���$��
���A�u�ZÝ�:c޴@�uޘ���즫 �r��w#�w[F���_�<����A�w"�a~���;o���e�{q�|2�������z\����A%�8��!�8oGl����+y�͙L���(�M}����p�a�f��d�[9E�,�Y9�M]�c��e���n&�9���diRg_��
5�n~�y����t�ݐ�Qg�a�ϧ�{���Am!k�s|yE���mj��P-j��X���oe43�E�6�=z��><=��.Q:��&�9�w��	��X[c��� M�<0��#Gܮ�{�vӞ=^��/�v/��9��;�	�*Η�;����kvj�"�G�J�i*�6�J+
<9F�li�t��ܑ-��E��v�M �]k|�M�q	N����<�s�ir0���;���`��䇏;H��XYED-�t;�πɅc(��������Ú�|����~T�]w��c:r�Nԯs+�dXA�Rt�	�v��6v*��u)=�R��/���$R�]X�;�¯]�))�z�U�^��ޒ� hғ.q���6�;�D�A��x.*��\9�l�5��X+S;� 2+�[�O�2�����ҟr���i��b8�l�͌V���zŔ�Y8GL��v�I4� #�G��H�@g�T�/VUy(���d�Q�K=� 1=���������ȳr�1OF�E�*Xk��fn��ۢͿ�l�.��~؟hQsQqP�r�����NQ�3�O�m�1T>��1��G'���h��
�~��"=���-׻g���A��R��{�}����� e���_��>����H�R�%8��ܞ:�fĂ��ɠVλk%G�vw��U(����nw��s���d5�.9��5|�h,���@5��ޚzqg`�n��6<�;��o�a�O��A�p���~��tK��,�3R�VQ%�qj����UF'4�e�yo	b���}X���h.��B����[��^W���m�����gκ?)R��Џ�_.Z$��ò���o�{.�h/���77��f�/e0���H�!t-�[������m<���~!��p�M��U����^&���}�O/�&(*���]����@��X�T���6��C��L�Pn��2�����_]Rf't]��	q�'�|� �/����@�_�|��^|�=��n�4����z�O���]�|���*2� ��y*�~U����ݟ�7PJ"`��z�p1qmZ0Jj����2 �co�ͦ=~� G\�h�9R�f[rY^cG�4�j���1%+�ĸ#X���FR�@����O�5��K����mzRf!�=�\g��ynC�><"}?J�����ʴ����]K��˔�5���l���@{L&���]ۡ-�B�"#y�Y�s?,J�R�]�͂����S�����`D�������34�h)����h�/�Eb��n�,�����/�U'��Ko�Y����qK���c����"��ax6z���|Z?�s��7����F�����H*���Sz�b�u��p[,a�����&�Em���`�hm��@{�(��f��s�3���A��K_�l^�$8W��<j��r�qI��k�]ǀ�)hue���Q��_��Sك�� �"*A�EX�Z�����W��Pֿ�FD�ɍ Gb4ʾ�v�]c��4χ�$�2:%g�4׉}rr���nB�,�~��:c���о!��v=@�'�� ����P�xe/>��5�+D/��o�D�'ۄ�$s%DR4�:������l���Ԗ�-:�}��iI��d���"�-�-O6����4�%ö�a�=R#×������-��䮊�H�Y����F؟63C�
�sFh��7�[��]��#dD��;�� �����-���{|�ݧ)W/^��$��U�[2�e=7�gQ%��7��Mט��͎97�L�q@3�^���d�*^�+�w���F������p�,�O�gmr�_�A�"e��*e\=C��X�Q��P���#G��xZ�V��6b�i���'�d��'\жI���l�@�=֒-դG�S�r���B1��6��U��`�����Q��d�\A���	�ʱmJ��q:�W�W���i�CǤ%wP���q��l��,��q,g�X*�Myz�ȪL��od��h1���p�։1�2�b�?M�E��PT+��ku�oՒ#ŗj�!��?�6�~pR�^JV�;B�(�O(�e���K�m��̢KЇ*"�yU�,,EkI�V����~!��u��Պ��jE�}el����Q�v���~��=S�0�ˢ��(T�?:>h�(c�y�=Hr䈷_�ج����V����
��xu��J)X0��/�f��k�@�<5���d��/|�����h~����e^�@���;B�󝟜�#B�{H�pǩ��6�'?t��M�Ɍ���7l�U�t�Jc�����Wx��hޗ4jQ�j!��*6���k����(�U�rt��98��|d�m �obȉ�V h�C6P��#Eq*}�a�v��!%X�6�7��� L���٢��z7��&��ܱ���	����_��݀�d|���m���bYQ����J��5i@�H�I��D>�E<g�3�it���Я��P��g���zL.��P[KT�f�;F�@/�0 ��js�Ӯ�գ;j�=����o�'I�I�6�Mu?��}]��������Җ�q#�L�煮�ȗ�R��ՠ���PoO�Y+ם8��y�/�sg�O�#��҇B�������C�v1d��
Q�Y:ѣ�D8�HIuz�Y�u�۷[=����C������T���0�ؐ+�\����'%!��Āyl>$�9j��N�����X{����zZy��'�-S�6�0��H,r{7R�p�(a˷ZI��k%~�� �|̷�����.�V���p�q
��J�S	�Lg�/aHd�l�9���z�=�a*��*�M���"���s|�G��Sx���������Յ �_{�=r�t1}�,]k�\<��hHND�f�ш�:�[�����d��u׷O�l��<N���O�?�vV�j�9"\���v�3_�L��V��h�g/��R��۶u��pB\���m�P�,��M_'h�����>�����/mjx�a�]�s��$�T�QZ17���J��2�bx�Zo4�za@i)^��5%�|��L�Imb|�Ŷ��IU�wj������4���4�/���͉�~e�<�v��#������94�%��-'qwn}U�J�h<����ܹ}���V������2~ux�TB2+�"��̏� ]�d@!G�|��:�L��+�x���'*_Y�����$�b}� ?���:O�/��=�'����c(�Z��Z��`�!(�;2n��2��;`��H�#��U��]?O��^C�N;mFa����m��E�o@��6���o��xr�i��f���5^4����}ᎎ$*�$2�c*�y�/���`ɦ�'��mp������ĲX��;���4N�򜔻
�+�>��E�ˏ��b��%:�Bz`�4��ulx���k*'�~��ݫ��p^i\}pR/۳�h6�6�!�(�����Z���K�9������9�}yH��GPA����
g!���<�::�ݒ΂(U�8"���T�q�=_J�}w�P����e�g��c�ʙ*f/M��޸E��,��M�͕��9�������?��dS�|���!�Y:��F���r�|�]xg�<����y���>����{=$��ͣ�? �
$�AC����/�>o�sd�����,��ŝO���M�F���O�Җdz�c�u����J��W�w.���a3C5茡u�+��k����M�c�%.B�)��]RW���3'@=`��D.�X_�졡m�sϞ}�iMq%HܡM6�W5�1ʱ6��F�MG���^�Ϣ���3Cni��Ox�ć��'��!)Pz鄎,Y]���?�r�f������� uS�L���"i.c\#�iꞃ���]��/1erH��J1�-S�-|׎�pB�𚚺���[�8�n�dHK;��$��Q�+$b���M�N���4V�����V���RÛg�f0Y��&��d��1s�?�~���G������It��6C�Q*k����r��C��]�����W6e8�z%�v����N��>ުG�L���S����ƨ��iK�!���u�^�~u��3S�蓼D2�]�c��^����)Jts�IY��[����[r#��4�R�;��p�1����KTǥ�Dy��V|+�J�R�Ԛ�t�� T
F�*A��e��:]�=Cv��k�~� j$!2+�~����`����1������x��P��!�ִ���{�|�Z�5����$�z��+���٘��ux��3&�W��.7�u�~�6��m���*'�n� D;c��l`�.g�=�g�I���:����T�:F�Q�ܟ���Ī�	t�|���g��nx��6�y	Y*���p���e��T��@�>��x�v_	�l�8��P��~d�fZ��h-�k�TMW�-� �/��cW�XД'����P�w�_�t�( !%�&�\��R0"�X�p PÔ�����V�O��P{���3�u������!��`��+{�2_�t���fiF2uI��,�f��Q��UK��x}d�F��h��^VG�2��W��a^a[�(	H�&݂��N�An�
�����9'(�^�o�2? �-~�s��ಐu�fJe��I�75fu-
���Z�"I/�+�'�����5�����N6��"j��)X��	��ᬈ�ג��{Ɂwr���HP(ʓ��x��8[�-�0$��_����Qғ���5��mˬ��e�hH?���4s �d�y{2�I��(1�T3W�M�;�/QQn�dn������#��*f���ضD97Y��Z�E�"c+�=N����x�sh2�q�%�cZ�h��0_3G���ŤjP���4����[�l���QN�UǢ�!�X�m�݋�i3�T��.LAW����K����v��D���h�G�e��Unp�|�5'��������h���)2RS�)3xG�'���k�E��Q\x�����9������4\<��邏 ����&Y��)�ض(�Q [^����E5xz
I&*[v�%Åz�~�����U�WvH�@2�%*�?�!�2R��8�V`���L�*�@�9�e����<�ETT�GB,=@ӎ4ۈV�ں�	�e�{�-��Nm$32z`������e7�t���kdV�KH�~KЛm���@<�,�8Ձ�.0Ͷ�S>�]����p�<����m�㕇vu�W��,��E�J��`��|��oeo��
� &/�*�
_�Z	��Z�����e�^W����3��qc=�{��Jŋ�K���I\��+�'�B��c���@K��nkV��A�Td�������$s��nzy�Psl�[e�f�;mΨ����7����T���$�r�?I�p���$�<Qg��A�O#��>�A�r;�?,�V8���h�C���Z$$ˢ� ��J{?x����}��"���KE�=
R5�9xJ���66�^l!���!{MSsKG/xB搮��(�Ҩ���HC�ԇU��,�.��m�o�U*�+`��j�<��0k�9�']w�О��SK"f���{�����R����^���Kڒ'#Xwu��H�>^_������p�m�>wJ��R�����[�܉��q�lx)��k��v{���u��cD
d��|�>�G��?�hd���@�}X`��F��X�״��z܂�����^�rY
�6�w��x����Z�;�q6�hlr�b��7�Lhҋei����o��=�	��e�h��Ft�<y��%�H�fQe��M���9�7�rY��Z=�v's�t�$��t�U,*��~֮��տ>«6��U:��}�ˁj���j�_�c�E�*]]�N�;�hӜ�_�;�/=s�_�U�RC[��1q^Mݽ8�x`��hcj��D�E�z��U҆��Z����d펳td���^'+<�Y�1M�B�KH��ӧZ?��`�~}��)'��HlةW�nV�̏��L[z9{�; ӕ]뎵AV��݂�x�9��A�UZ���~0/z�hU+'��h7�	D�;�����ij����<��;�1u�1��oN�*�V�-�X�����N���V�)?����Ε���2_���T����oP�e��>&h��6RD���L�ys J�����Ls���a�b�F��ʺ@`���E����f�ϥM@ ��8Y��o������,$_��Τ&�11|@}�)ɫJ���Sh�Y'�,��#���Cz�PJ�n��Ш�~��Hͪ{��|Pg��wI�TJzE��߮���9�4�AB���Q`�".�S�;×��ns-�q�P��3�F{��W���6�b(=פ�-����I�N���D��"�Hk �"?Z�H�뉿ܡ��3G������A��fhx
+1,*3���^W{I[
�T e�O�3��vҹ�$j^��ؒ�g�(���
sY'V�v�h}ZU�-��^9�^uT����@�5�/ܼ�|���0�B�ܿ�ǲ�?oI�(�Sp��9��Y�Եh�����r�Թ�ա�mKH�%KEU<�l�3��d����`�J s��Ɗܰ��^ݗP�m"�w��4������; 3����:��g��o��A��rE:*
�o�A�i�Lݫ`_b�$;�t���q�F.��r;0�25���;\���C'���~ʶ=h�v=?�%}��	�7�ֵ֢p������SI�WQXx�����K];�{�tTx��4��S&%�?y]� I�9�淵?���pV׼
������feS��A�RW�A�Z�Ž��f��t��c�|^�sCm���3��}'�[��Ú����m�=�~���_��8��O��Ja�R�S�.����
F��W�A����ҹL�(�z�=��/��ԾG{�*�E��QxC�A���bQ���n�ݤ�ܼы �ؕ3�2�b'gi��Q�"fz�/8�A�US�����˘��c'g|�K���<V�����<jMBDa b�|��gnrvP�|Q�7S�paK��yU�^X2YE�bӮB��Y��f���)��f��@Z����;�FV�/��aW�GG�%�ϲvaAQ��S%]J��O�_�_�_L��?���%x>�q�Y�sciwp�<6ϧ;Οx��}���S&/�B,*Eô.���oò1)�1�����
�� ݓύ6��h�h� 7�OE^x���>m����Dvk�;�O�U��}���^ӣgM6�O��͙�֯�?�/���Q��W��D��4�ݹ6�ʝΓ
�Z���JF����_��r�VR�Y7��1���s��o�p��(�Dji �rHћ?�s����_���}avJKy;�b�קӃfe�b�Y=�k*��'>1~Uro}�[e	�����F��Ϳ�L���/�1s)��3�
�}�e����5��Y��Q�0+��n1�w����~{j|�� 1ɔ��th�T���|}��~�U�Z�]'�u	�U�[�-���Cȕ��x{M?Lg�����(B���{x��ܱG��� �U� J�����I^[�/w�� �m�j4���!�7��u׆t���6�y�o�������g�x�vt�i�^�^�޲Q�c����#H� � �=,��Ѡ�Q�+�,����F���b�4�l�����7���uy�z��͟������ݠ�hH��J�л��J�RwR7S�����2��etq�hӈ��;ʦ��ISbYP���-������vۥ�~��e�Rb
G�wF�����L�n����h�e1�쵻�B��9�;�Y��+���5A��D��+�^z�[����W&Ax߱�-�o�ظoT䌡v�����!�+쮙	p�����f������u�;�F�F�S�X��PŘ���E�� �>m�'=�e���Vg~�V���׿�\Yd�U^�x���:���G�;`ᰁ]�Kh�1����%���	�k�M��?"�_�#�I�`���́	�>\h|��mlь��w~x���b���+�͛����Q}�Z�/���V::�98�V�/��
M�e��BJ��:�{�wA�#��(�F�~#�F5;8UT��9���lA���������;�]7O�J������"��	��2C���Ho�)�� f, ,,<,�����M�!��n�F�ƮV"�<0g��t�k&�Q�W3Q3��y,?&�䄬�%�56G�w0�E�{��Y�?���$���:(�rm�8�\��ca|_�¬��J�~r�)]Q� �V����0��ϫTw�!]�nfoq\K�V1������d����۱���]uY�+�5�u�6��\O�>\���bw�ɿUҦ˷X8SsG��q#a�X�	aHZ�b��+e�����.^��T �f5�=�
���r��#���@EvA@7�]�O�&���S0�z�D�#�8���/�X{��}��x�w����մ.t�')�Y�3myO/|dO�s�S��KΜ	�V{U���o���U�vX��U�ZVF���հFϚ�?����$!�$�.QUC�>�gl~yR���9�vZ`�Ba�*=��͋��(+⬙�B*/�pvYX�������}v;�в��3��*T1H!k��,'�%n�d��r��k++Dv��AM:��I�b�FJ���*�F��s�p@w�o�'�����r��bۥ��YY����Y����Sf�<H�}vD��+�$�,�6A�c��87�#8�r�\Ŷ���\���S���XJ��>��L:KK�\�v~��C'tE����`�H���)~�@1M%�P�	'Q�Q�Q�rUZ�\���������J/����"|���uhs3���j�g	����'ɤ��8����_�MH��D-��2+�c)�NDёO30Έ��nW��'�3�Iti��Moe�VwyRHca�3�����	A�eJ���np[8��s���)Եr�RV`��щp� Ta�o��Y�:��,۩��P�����	�)�{K�5W��3����Au�	n]�=Mx���b�~U�}@+�����þ�{U{i*�0w˹']�֌�Y�J�+H̟)��C}P�H_��f��2#�̮٧��p��tNT�+��B�VH1C�3|?gaQ��#G����@�<Di"���?��ڎ���|�Η�Ncu���^KBP'�.�l�0�ɂ�0c��i�f��@]/q���d���!W��W�!@
��t�����p6�#��M�ؾ*��Y�r�1QYp*��VTCu���ҭ��{�ɲ͋�XٯtiC���KQ*�X��M�м�G\�ܯ�1z�8R�3$���{'�\o>������6���������"��mc&��W(9[q=����>� s����P�;#��^m�S�o�(A�����^U1��j9�~�;=�%�l�>�ŨА�i��D49�(�5�����!���C^(�.z���iGG�`�AN+Q|������X����N	�r�E=��q�x���$�is�Ċ�ݢs���а� �d�P�Dvg!Up��6t'���_-j��=��E�m�ŵi	Z��E�z[�[�Y�Yס<2Y6R�5�\���f�Ь;�t��T?�u������-����t\���<)4Yi���w1�wo��#�j�6�5������i����N1o2�H��l-���K~��K�	�wp�z��ʶ��:����z��K�|޲;{��b��ͷr)+���ؽ,�˫%����i,���YS\��b}t���*���ɢ���ґ�E�&�����򊒹��\�� ��<Y6�;���J�����D�	W_��2OXs����� 3�^Ҩ�\L)�RwR��i|���kLI־�!skr�n�� �UMz%\��0�~\O��(s_��w��e�N���=�B�w m'L��>Q7+��g/�O9h��pI�.�;���s�[� ���Iy+K���#s��6k�o�<A�#�QJ }��+,!��d>�'Iƭ<�n�K�5U��_��3�o���&�q=�峘���up	5*4b-R�+��b/��G�O�O���Ok�W�J�� �QR$Z3�n7rٽ3g�xg�p4j}+�� %��{%��E� �:A�M�^]Bd�3U��{DnD��	+U����4F-N��So��p������g!�i��2O S��d��T�m¢���g]%�G��[l���1w���	��5qW�bl�ƥ!ɯ�͋��Xt]>�Y�N�п�[��_�'�>���7��<� �R��4�̮�К�W�h�_�g��a������T��3][��5m��ƀ8���"����C7Is8p�k[�/?��3=K:�ap�p0���nۿ�s 1=���m���f�0�Ɇ�Fb��sp���׵��mr[%�yH�-������	����%���u��q���I:�fh��н�P��f�I6�ʱ�l���V�,h�@��T�B�4��d��>�In�����+�Ύ��\=A=�5��2�F��[5�� ���G��J��Hp�1��瘗&�#������`L�w�jo"Pc�kym�P�ݛ�*w�й[ݒ����2�r0q�|���E�|�f"�=�9�LK�1����'g8�����KF�p��?�[ǡ����+�
A� .l9��Ϣ1�O�J�tϮ9�hg-|�C���42zЩ�O���zmDEL*g?C�}$�{�E8U�b5���CE���t�;g�G�t��wG"��-*�/g������N��ڑ����`�y���#7?����e��)N�,�C��>���0ݯ�RH(�:�����mb�~��H�gr�`�M�b��d�,��7VO�Xk�,�~a���5j9���<�7�_-g(`���#������Z3��4A�)K>��;k���[�;�R�~g3g���K�`E}���O����:�w� b(U��7L�b��
{��)�c��pU4��y��1{�Ğ�.-@M��	�	�����D����#�r��\��d�������M���[��zn���|���,UV�K� �S���|�h��A����ŖQ}�O��5��M�>�����D{����*ш��4&�}T�+Z9A��S�3O���� N3փ�-�7��e�\6�W�[:�e)�!�'��Cv��V4� D݂?��7f�xDb�J�7���~�_*���2 �ы!v�B�C�b���Il�U�|�.�ڭW�� #)��X����8-�ׂ��k��J,���_Q�k�ﺟsG,�S6D,N��Rؾe_�+�[��OIGl�ǀ��)�A�9�a"g�uG���y�8n��ō��$](����k��O�,F{�R_�t��6�b2{�M�y��^2h�C���K�[�������nTK:P�R}��E�����6���Fв����cҕ|����;I�O���5�����d/Ư���K�p��gEnv��A�m��N��^����2w
�N2����aH'��Ӯ�A�����c�$�`�_J�˵�j����v�!����؆t$7�U���)6��	A#���Hv���t���c�=c�4y	��є��HWp9α]��'(5G�S�##��뺧�	a�\'-N�y�F�m�q��r�qM��e:5+g����R)�I�楛��6?Z��!N�V-��z���Y�/�.�NK�ZJ�!I7�Ö9p��(`�e�.��1�G�;�����돿5� wߢ��u2�}�����������$/�9
]��DPҏp"��'SM�c���hI�酃�w 2llY�4m �<�h*�}�^��z�t~�!�&��dwÝ8o�3�Ji[�E4��B��_��������$Pw�=�YOZ��>��{�h-0弉�����iβ�O�a�!�W��x4��om2�6P��ʿ�R$���y�Nds�L���R�P��f�s����9o��q9�u��;�zM*�b�(���i��d{N晉��ė�#9�F�⾳8�	}����Km����Lb����`��0�(�91Y$^ �cC$ղ�D�Ձ�!�z�Ԟ�5�@baf���K$��s,�|������U���f���!~3:|��?�T�ˍɼ$�*�v�@ϣ6CmZǦ�l�<���J��C�f�&mWŊҤP�>EI>g��1�k��4c��@�Z\a])ծP�a_D�~5�-�-󝉁���-�BI�*Բݧ�OʎP�T���Ƽ;��8o��(�O�D ���auB�#1���.�ǀ[mc���W-m9&-�0�C	/��yu�ׯ�Ț�zR��I�E��Ζ���f�Iױ��F 2�_ZA�Nł��i�atf��ZUn����|SG�*��j8��9��e�����qb�����J�хh��Cց�ʾ��w�J2�P��%�-��"<�i�P�^��[eZ�v��.��R��*��$S��;��BPA�e��7f��j�6Ƀ$	���/=J3�n�̺�)���d@�+ǖ�U�j]"�f�ѾF�%O��.X���tIM��P�u��`��x_|�)r%�F�e≀]o(���>�$��4:�=$r�ǃMg�m�����)�������YM�ޯ����]��?l~B�{mU	�� ����+��f8[�4�*��"�V�D)~a:�5�&����8��N�#��%s�1q�T�g�._0˸�+G��߱GX4��tm9�+H���TD�r�]TH���%������QZ����p�p�q��r��3���r�]�W,.3\!���*+����I�`U�������p�:%�cƸv��>��KD��`�0",��w{�L���#���������:��n��Ul�n:�FmΛd�??�������`��<��
;�Uhdf��F9�H����[��o��ĝ��cl�X$DW����Q.L#x�����gl�N-�7�No�.?�pW��}��2�Ĺ44<��8���Ǯ�d[���(~ù�g-�~� [��S�e`�gU���f���sI��ouR'���D�ݗr�f7�<����$/ZN�7����^[�b�H,��>��{���8�Kt��oD�P�'�<����cc��8�#�����E1G����1J���D�PmGV4���0�~x���|�{��!\⹭�����=�?e���D����rr� �'���w6�?TB5*�z�A���M?�Ԥ9��uF#�{n}�������V���k�Q��g�������Th�%�e��WȋC*�P؆&����8���$�]���c?�Oc�(+��id�y!�pR��F6G�����R?Qv܁]����j-�,���'l�>aDj7�Ϊ(�6O�P�2�5�_d�Ξ���';9Π�܃zއ*�Ö�k��0ک97����]�	�8H�漆J
��2�If�a���zg��TT�<Ҽ�"�[c���-���G��3�g�����M1�b��_�|�/u����9���K�n�1E�ߴU�4{�8n�Fg۷��hYO�v��z��Ed�(�o9�l���ym;�������L�3�8oG�#������1�"��Q�͋l*�?�$.����
\�Y��Q,�Rp��-�������+�q���u:?�0T�6����
�r,N��X�TϨ�¾�'$e�P�
�l�����������U?m&z�Jb�bW�N�1��G�Ɏ��(S��<�� 7� Z:r����R1��Lvq�0�U(ч�b�U�N�*m}3:�[�F�v�`�l�c/^�?�eT\M�.xh��w� �qOp�F���5�n!���,X�4A���@��!	��~�w�̼wf��;kn�^g�:��]����]U?�쇾̩ߺzk;��j|y?$j�܄-U'y�*P)0b�Ȧ9��,5��p����5)�v�����ʩ�Q_eo����Ʀ_D�f��"+����5��H��H���;��o���zB�,�.U��}�4<clcq���<t o��@��}[���t!?�����+�F��&������w�#^%>�l�uޖ����ES�,�,Kv{��M�jӓ7UPH��vNi���k��u8���UvK����ohM��Ẃ>U`g�~|?����| ��2��A{�m�DvѠ��^CqG�sE��΃Έ��w�XB��Ɯ-k퓵*�N�:V��o���ݓ}yQ93ɶ�k:�&�:g��Ÿ�)��c���yۯ��]Σ��+�dY=��<c�:Y$M����%��aU�'l�Z8����I����Y<��?DR}���)���Ò�y�҄����`���0,��ɖ�%��ç; �@5�yK��x#·:�s�u=��G�?{��"|J��O���9��_;�Y��i�B��y��E٫.�vk�u���-o�8W����� G����'�S(�66G1�p�S��
�/lj ���1�B�~�~-,O�QH��~<���(�i�=��NWW��R� ���_(	WC(��e�AQ��y�yb\�����1��~Cz&{'}���⟹�j2�\�v�Ќ3�A��I����ѧ����(m^�]��ݲ����-x��/�G�s��IW�i���(^pH�%�P�����ړ��� @����� ��Z��m��aJ�뵦&UL�`����'���2d�G��C'Fv����8�3"�4%H�_��)�G^��c� ����6��!z2�,��8MO�AR��(��3�Lxp`O�G�K���JSp��x̱�Lj���d35JIi^�T�!�>�sc��#
I���Ȫ�;������s4Xv}P�C�����i����}�aNI\E�}+�2A�=a��U�11u�-����ၠ������f9jql���r��I�O�	�f��A�K+4٘��+����sf�a	���T_0���&��YU��|T�Gh"t��oϐ��?�l�����M�ILM��5�0��:>���Kj�"B��b��NDIN{���M),7r8�Knܬ�?(&H"GAg�hw��7m!?�	���r�Z�L�S����1Iu:�CFJ�+s��2I�b.�|�D���j�\^�"��醦d��`����:��D��"�a���q"Z���6�H�
�yѹO�e�i�׺�=�c���P�p�$�㖐�^�ݫ�����:�FbK��^��}��)��&�i�
Y�;��2��Z{*�R���ℕC��㞤��5�-M�_1�~�6�ݗM��&f��
��p�����$���U{�اJ
� �����x~[�k�(s��Ќ��I�A�L�̐G_������	�	�])��h�9�w�5�~��$��oԸc�5���/x�3��(@y�z
�#s�5�F�lي7a�bB�g�B��XϲХ
�FQ_r��PV�$�����^�:�Ľ�l��W������n(�t"�x�^�"�!����/��d�V��2q�&�?wg,���Y��@�V�fjύe��+�(�Z8�SVka��c�s���8Gt`�{{�PB��v���4���7��I>���br�
�J6I�hgh�GJ��f�kq,n5Ֆ� �G�N
%��R	Ŧ�P��*WO�õƑj Cn��O�K6�@��h�piFT�X?��D9����z־�l�6q�P*F?ޅzU8/O�e*neIHdU��W��lVY]�Ÿ����Rf�4c���b��aq��h��C�x�
Xt����e������>ᙲ[��+������������N&Lz���fBbѹd�ǔ������I�R.�g���m��:GV��kC�:/�ڇm�"�J����*f�K�zdwV.���.^H������#m��̎W�xV�2��*vÛ�
�d����s��7���sr�DO�_��G��j�2��܇'�֛���/�쭭jru�-�_�{8(���*ɥ���� 	z����!��ާ�oc���mk9`�r��xc/�O�3�����Rb�h��5�A4y�=u�j�e�4/q���������?����
Y�n�w1bniYtUڥ�!���T0#� ���6�ڸBB1�ďe�\��0����Ģr0(7F4ۛ���_Z��E̲�5y�ٔ��3�	�th#,Д@��N�S�d�����ßad���S]���utC�h�e�!Y�C�"��3f
+��1\�l5,�^d�ͮL���nNGA[�M9�W���!�cǸR�c�O���,�֥��QXuM��l3jzu]J��C�.u�QO|N��N�Yғ�$$��FZ�@�^�$�H<S	n"�"8����(^����U�-v ��O�Sѯʄ���}�W𞃢�\	��
�²+�����"������������Uz�Q�T!,/��1�qޗ��������F�^�nA�f>���ϩ�D����9���R���Z��儉̖^ ż	5^;d�n���S?[�]�k,2�26Mn�:��^���V�\���RU�;���\���9���[��_��/�~��;?С�K���^�.������n�nt*�ʨ��u�]�I��M��ι����zemx��z�]n�A#�����H�AwO���z:O��@!�ٵ��I�\�E
�+JB�Y�nP'Y��{Nq�N�SG5C~��Iy_�/�b/)���³Z��I�������A�Z�2�{�9WI&\x0��$7«�L&ho�e���姎��i�1oH_��8�����7?� �^��]�ԍV;��J���%��&"~,R����p�A&��-W�� �����5�p�V���9��d��������bD�+(�D5r�̥X	��ʤ���b�qr��F�mɶ"� 1TGd�3�w|uJ)z���7m�[uyz����Lz���5���e���:�P`slO>,��$.}�+�~�����/�~:m14�0Ѝ^L/�/(_hV\DV]� ͗��n2�9L�n�C��R��~���]��+�Ky��?��cU��e���)�$%�8Z��y7N���������u�±��W3�KVa�sŒ�?!ݑw�_Ec7A�/bY���A�L�m@r.�8+��Qщ��X�E(�S�hUm�pC�ѩK@;k|�ejj}{��'��I��`R�m�/X���Me�D��lۗ�.s���E�k������I�s�<��^�/���v˒�oD�e���e�k�Oa#��Rx��Kn�u�|w�z�1��Ͻ̵k��FY�YE��R�Iu�όG�l+�Cy����(��Ⱥ~�8@<�ݝ��>)7Y��$�ރs?AoƳC��0X�$?����F�Cȡ�G<��bG�5�͋Q�}�́���G�E �~ؓ=�"/�_vb;%����Q��䍈��c!��;B��R�ڃv���/���U�m[t�u�Q��0M����lP:�Z����XC^w=r�H�Y��ٮ�ŀˑG�Q�?p����w�4_��ӑ	����c8������L�@�/'����^N_�o
��2��s��k�z�?Hl�Zjd�c��A���H�|"�AB�k!��%q������\���Ւ�]��r�9J.<�`����=t���TQӶ(��\pcL���C���kVЛ��l��H��*a����z��{��Sk¿*�mh�S�J�J�⮶�j~8��٪�᮷�� ���#���FP ��a���D4Rٺ��̘a�,���F)A�a�w���E+-�Ƒ@"�[:�E��.>��\C?Qa��d�.9�%eR�|N`~�u(�a��S<j�f2��v���#�0���/�@}����~k��#z*�&���+��`�H^��R�5׆��2���s�,ߒc�nTZjѼ�e#�~�����5��Œ^�G���t���l�'ۂ��LP^Q#S�:���Y����kmƌgV�A]'K͙�Ʒʵt󾐾�Bz�������GK`�t�QM����7�&�.�ג���s�I�z�QA��quZg��k����^c�Br�g�Ʌc����-�9���?l�k��S���Q�8��݌<������_�(�>[��Ȯ���:�����_격	�QQ���N)�ϛ/�2<��$��9Ƨ�+/����,.*B����j�Y^Ԧ���Z�10)�Hø}�A���pS �_�J�.��y4>J��������"=�`���ͮ����+��SB���R�
����+�
��W�\T��>�C�w�`&9�T�5y��/r0��5��mvE�\�a�; ��Fosq���� ��afmŒ������2X@��8��r9Wt �Զ��.�PN����<����� �����x�K��5�ǵ6W�zɔv��_�f�<l�՛Rp�+V���Y�Hk�˧SȹDMS�膹"F7�0�"hu�o�`ت+9�yv�>A�	�dG
�=T �Խ;Ӻ�I\�
 �x�sOD&N�an>�C|�Kٸ����/b���ڿ�����^�S���M��]����PJ�c��/W�o�F�$����l/qx�yQ�`�j&'Z�MS�ւW�{K}(BM�� �������4�����G��b�'��q8F�8B�����	Uh���Th!�*`�3ny҇�G�.�js"��g2*�2��lK=3����A�"�&���m��TdL�K���]���zY�=�'��t7�9�~(#��uJʚ-�ׁxQ���2/��Q=�H�Jk�h�H�_��� s��e��*s��n<��<���u�k�v��F��n�{�Wc҈;M�&JwyP���Za�̎���H���@Y�2�ܶ[�Î$��]��6ӑ�*fV|<4��T�ݲ�
C�o�gH�k*^��f��F2�a��;�� ���x�����_�j���T��(�K�1����.a�C�hޙL�ay�mk����l"O��!yߙ2y��v���E�s,�}��"�`��y�Y@@��=�¯ڠ�
�^�hH���wC��I}���#��oc>��i=�R�����vA7Q?ԐVN�A齓��4�.;4xjQ��,�(.���}~�{�Z9|�������@�ZF�9|�w�ʿk��##%j�z�2/{�D���G
ٜa�g)��l8]b�-�]�(`}��E��Ɛ���>�T�(���,y���Oa�x?ND�4���ӾC���-M6d�|����W�w�CJdV4�J�s�u�M��1FR�D���gָN0�Nμ�������l ��j��OK8o+w���+AjR�c�]m0�E �h�-s�xiW��=EŽ��LA��ȑ�����'���v1�M!���.�z8(>�f'ͫ���G���6���U�S��o���ER#�k��A7������g�²������Y��2k���|��6������3;���l@�ܑ���D~X,4�#O��c�h�X)���1�ك�|4S�K�}d���<-p�=��}xgX���K�o�qP'\����D�gKAى6�F�\c"Z���w���;`U��W�~����/UR[I�o�W"V%��H�N�t�v�j��ȑ1��pV��E-�X�7ym�e�N6o_o!ܠ�a��gyu1Oo��s,�pr����s���˧�Z�?�	�z�ڟ�mg7|�葘0&!ϩ�����"��y�K!C�7���t�zI'2���dt�/.%hۡ�R��EI]Ʊ����x�Z7O�������<yV;�Zh�t��ڣ���4ք�+5I�>�i���b�%篳��V=�n��	�6��
�w@��75�[����	��nܶX��)�8��F`��+T�_��iwK !& ���'����'�u�.��_��^����6a��p�YSh}˃�E8��U=Q�f�����E�dOez�J�3v����!Eewj��*�Jw�4`*�Aa����QN�=Ŀ���:��-(�"�/�5"��M��� �Ġ�ӂ�i�*A��ocCYMq�l����J�V�&C���-�	���èH���Z�ӂZT @qU`����G
���=&�0m�t�c���7z��҂Ơ���~��р* �`v��3p��]����zޑ@��,���"0����c�@>�@?�K���LC��ߦ!E`C�{6��0���j����w��#���l��׿��Zͬ����C� ���G�I4&�R�I�ߺ���_��`Uȩ�7e�9#S1�x/�V�!�W0�>/��<����{
@�P��x�5s�.ܢr�7�֢w ��<u���?�s�Kg��� ���yOCͅ�� ��KnN���*� � ����B	��@��C/INA�o�ZD�+]�����D������1�y}i?⊝��4��0�ʿ]�c ��Fsp/�@	W�<���Z[��%��/4����1�F���G��4B�݀1F�8�k߫+�>v�?�ʸ` ��e�tm�sH=�"*���:{�ҏ�������k��"��y]�-[�c��hq@P�,��p�]��4�W�A�0@O�G`�!��������!��z#��&ϭ�OQ.��MR�(��L�S���M$.�H��R�/86�?.@�Ă,$8Mx�0���"�<)n�	��)#�g+�Q � И�K��� �G�f�s���qQٟ������}/��\Y����O���8�@�гe��sfp�v���y���9A�F!l\��Mq�+��8B2%ؿ�`CA�P�>] @@�m����Aa`a���տ��f(Q]�q@�X�A��7�s�2�TNz��e�t�x���ǁP�~R�Lտ� �  �� >	��� p��j�h� �������H  G��(H��`��B��OE���:�q/�p���C ��{n�b�O�ӵ�a��l�1�#�Pt�>K��/X8R����l�< �)�S�Zq�XyJ�%�DΛD|��o6��\ �� M���H0��P��JOKk������n��n�w� �?� @����!�����L��?�A@n5�.O 0���`�O��� Nc ��;�-
��_��?e����!�6|\��C�1z����펑�j� ܮ%F����(ŰR�-�8�M�f [��I��L�֊�\'x�)�{9���!0�́�A���5Fv�����3�~��2�*��:7*Ҏ���H�p��a;�m aۮӉ7Q;�Ǩ���S�#�qMl$�e���R �w�� E�yf�T�����ԗ'XL��= �I?
��F��A1���AmC�C�A#u�Mro@�{b��y���Y "zPa��\?��2�ܪ��s�Gܧ��H�1VV��? �� 
N�k, �\����*��`4�F���!`=�V�I��.I~�g�~ξh ��Y�2��	"���_��]B���Ep?ݳ<�`0��#�? ���@�A��k ΅��⢸��� ˒ �Jk������3e�Q�_7�Y7���bIB�'�*��/
S1qK�U:��yހv�`t�
|�5��@U��!�gy�`LW`)`1�g�1Y��?��+�-<�)�W��҈���2��G�o�{�Y���^��♚}���p���ٴ�Q�D�@�?�lq���������|���ON7��q`�p���j�z����&���|5[q=�(zv��t�4����0K^|�h��y�{.8)ki�roT�$�П02��� �@�ˇ��^)�u�!DB��l�Րzo�vݣ�M:�e�n����y4�����MA9����{�d�?���{��P�����gv��+�&J{^l�J�D��"����¹��-�\2t\!M#�S8OP3�u���2��xo��1�Ԧ�5L+���hP;Q���4r��D��x�o����K���{����!��w{�PyLv�4'�u�����I�;�N<n�P;��`����9�x��C*& �QJ��s����)Y��1�Z·��Yз�zyT�{�^�F��L=e[��I�m�T��*h�p�!�Æ��"&"t"x���DL.,�M��oP<I�C�'EF��6���hy"��ɕ�s�n�~�~�Or,��S�{D�a�`O�ㅟV^���D��Xd�����XvE��A�[&�tf	�>���t�N՞�����Ӌ���{�1�Q�YtZ�GT��g�<� �ڡlJ��Q���p*n�y>zƅ���Tj
�AWo�+��r��U�{mz`X^&�)=�GMn19�%�G�V�$v���tX�Bd�U)!�� �5��h�c����}k�_0͋xj����Nu��:�a�wJ��<u��E��i��M2v�ި�/v_����]�Y�H_fo�!�$�!)/[Mb㟜��S�]�	z$�wD��>�^��v�ܺ�-���*K6j)����	��pӆ.%Z�d�̾	z����ѷ��b��r�J�[��M�L�,��F��M�&��fc�^8�d)�~�Z��В��q@07\�ʼ�q��C�a||�k������h�u�V���v����`�L�W�L�U�b=�L�rF�]�v�Č�������H̤��aW	����� Nݱ��ʦ��^�5䖘��=�)�϶u��l�PD���٪LD9�E�װmv�Q$c"��K[�Pn��t�¯��;�0��>���[�D�*��j��h3�,	`-%�������P�uGF�O��-�Ep�O�iQc``"7��R��M�Ǡ��^|<Kj9�M�-C���/��ʖ��δ}����8�8MH�Һ5e�̔}c�:���M�ۭ����Dd���Q��$��p����I�O8X�5ъ[r�՟��iuˍ���K� 4��ZD��sN������3�Lw���K��H�̢�<�#m��fr��iA���U[��w�$_�/�;` �h#��sݸ�0xϺ�2 �2Y�B��ql$%��"̼�O�鐣`���{����	d?�Ǡ�i�{O���(��T%�䣢�p��0} $7㹺�|WWV��3��.�QW$)�~� ȟ�{y$�ǆpDU�h��0�~�K�2X�ˋ����/(��x!��(����c\_ۦ�˜��L<�yi�Z�-2�п3s�#ڡE,��ن�7dF�y�0�l�~X46VH��;c+#�.Z�Jhǁ�w���;��S�:�
.F2�����Z��
���%K���9�m���wX��6�wUu��0��秙�~6�k�7J䋋F�S���X�(��������'���J��t�b%�*l�y���Ҋ�}6�%`������c�b<��E�N	_���&�����&('~���T�����Q�̅�Dc���㜘�!�"��ԍ�劋Ű�������$'��[��͂&����N���#j����d���-U��7MQ�RW�S�䋍�uo~����5.2D��H���n���'��PՕ�d2�ޫ楣s�q�W�+��FL����	�PԆ����V�^?�h�:!��L=��'�n��1��'�� 쳑��?1���&��m�_M��n���"u:�G�:���&e�8x=�Uc�E�(+5]�c��m��M���ލ�o���4����`�C�S�E��U-��Ţ�JG�����mlZվ͌�*(�$fޞ��[��sYn��AT|�ʒܵ�d1hP'��I�!�����G���SU���m�O^�4}��:/Bvy%\?J+&�+m�Q������c�cC��0�<�J������Qj�:�7��g�7rZB[]+�5�`U��>�`������zQ�6S����nd��>`�����V�T��=�(�;L<7f����4KeU����4���z�&�u��y( ���hn=$[mҋ�Z�q�p	�ٵ���ΊїN�^/��؞��sT�?�ӏ; ��%�i��Z�I��%ɿt����ى�ٲ�xQ�1Ō?����ec1�W�U�b�u�T��~�V��jFW|��7�e���삓��Z��ާ��L9��*�ҟc��5�u�������kN`҂�gDjЯ�D,:�B���O��j�E&;��iY�����.�x{x���G����[/�1-���iY�Ʈ��"q)��\Sӎ��^E'&u>�&R'�S��Wz04'<�q `;����YcH'W�K���`�='�biYTX�w�D���á��'lj��G��/Ց��_7G�ĚgO��~�V�ŝC�<���1�,a 7�v�H��z4�=5P����'�az�Q�D0і�3�Nx�bľP�n�/�1{>�d~�0aP��K)i
�q_�!��?#�H��t/�Տ~��#��Ս8�$�u��C(2%�,6d�4�W*���h=��0=D�A_nS,]��R��#�89���Ʃ�����ja�G�ۀ0�z��<�����A��|\)��0���?�~���bҚ'�����t�.�cMx' �����0�=cP�Rd�G"�yފ�조�,��罂�CڞiX�6u�eZ1/X'��0�-�����(��[�y~K���^���EP��&PSt>u�SQ%��ʲx�DE|]���
��4���´�~�J�?�
��y3.��}5lLh�t��J늬6�P�g��w��
x�[x8����c�3u��l��Vܗl��/�����a����_n�zz�<�tف��ɣ�f��%�wji��%PU g�y^wf/�\�a��5�`M���u戉��Ɠ�����Xs��g/=�9�(�?�G���~�� �Y�Z�1#��-�%�cBR��YB�)��v�9�c����ǈ�(��JtG�{^�����Qhf����C�}rC>d0��W},������A��s����'�ϾNu4��w����q(�T#:ё���$��O�����r|w��z�M�`;l1�:m"z^���C3>�O{ɪ��q�moz��
�>����xM����1i���[��*��/����h	���d�����H7�Tg^����;�ADͬ@���&��t"\yP�dӡ�%�I
�ۗ��V]��1��E���v�ޣah���c����,L�N���Oi���%�����/�]�����O�A�ލ�2��׀��0a�B�a�q��f�������g_�^m>WM]L~�N:�].�Y�p�Q>6���+t�����n��&G����c�%�!��H�zK��q�`�M\��o6M��ǖ����\���> tQ���KS�'K���|ն����k@[xE�z�GU��q�oF.Z7�-�U-�Dhz�M,�]V�FB90?H�,M0;���>�D�h�iY���"~�/���1�:���by������`B�̣��k��x���J%���M�/��b�~,R�Nq Dv�^xqS.�G��z�f���U��}Շ��<�5����18��=�����f2�C)��OY�c8=�Ic�A�����亗X�S��%�U�O���4�[�R�s��5��7|Y�ɥY�Jr`.u�n�M��O[(��v+r���ľב{A&�@�a�
!V�Ud��)4�����^�tH��+��w��X��C���q�:=�{���C�V�-�oم��B&,��GjE�A{����Hs�9�^��&������/G�>���d|#�Cm��L�٠c�	�����[M˗��o9���b��i����w�X
<,������,WZ�Z�̑���y<�B�P�&QE��"%f���k�e���|��'y~�E�躣��C�Y��j����m`�[��J%-Q�C8lC�	G�;$������f*��*���%ٟ��pW��˫�W������&������4b�`Q(K��f�؆(�� ?��;�x�5��E=y�]O����|}8P�&A͎XW�_����F[�x�D�	N��� O��pX$ǉx��ۇ��Y}A��hVxd���$%y�������<-�'.٪�5")p�y1Y?ޜ
�څc��c9ͧ����)��K<�ܿ��4��h�Rlag� ����8�d� W'����_�rJK�"c0=?+��7����rr8"��@T���)�(NN����ԒH��yD.{��?Sx��;�-̮6!�-��"jm�<��+d廾(��9��}a;��~��z!�+����܌;@�<�����`���}q�Ο=v�Ů(˱I�� ����}��g���M��L�㔔�7yy�w�^��p!5��U׎���֬Vd�f���L���`���?�%���ؓ�_�=�sɻ�8�~�� B��B鄧�o��£�Fe���zH��SD+�1!d�9���C�G�ӿy1cl����Z?�B�M��	@��Vk��jfv����*���U[H����2���B򑤞�����4�?%U���"J�5�$����И6�^��Z<�ۘ4�� U��Δy{�x5p*XtT5-��솗&������8�W4Rs������ia��C��/	�![��|rӓ�zO��^���N8|���e�9>i��F���
�����e#�
}��ER	صL�7_iob��J��a�{9w�T����,��C��=Egu:���^7{l���(`��Y��K7�`���L�_�ע���-�Ҳ���2iZ�̖�	,�ޝ�M�	|+2��,�ab�S�����?�@$�Z��&b�YM���p�bCLEoo`UQ�[3y�;B�G�egGX�"Y�����]1̙`���/ �˃!�1�9GL���P��r͌v��u�?9�79���3)�1�JO�i����o�|�D=��l�P8�1��gݱ�;~q�f\�
�x���'�z�5��?�n��^N#￉|w�۪�4�ؙ]����D����w�iC�������E�֨.q�r��nI�z�I�L@�4*�3zՖy��If^�7���?��C뎹�@����UXs�J�PT�[O�}^r=a�m[:��4��D�r����%�*�.�c00���ނ���9=J���pt���);(�~�X�9��u�*�vU�M�{�*;��\�R3<�׳ ��N�Ӽ*��sd/�F��]����7���;;9I�;��tt-��>z��U����n-z�E�)}h,��ˆ����b��f�]k��O�����ܕ�q�/�C~]�w彞�;C����\�%@5�x]��ĨΎ�j��Ǘ1ӆ��SM���|�Y&�ܚMz�.,�)�+�gUx�������K���D�s꭛�=_�9�\SS�q����o5?7�͝ꥧ&�����Қ.^	�O�]��~ɂ~��@�KV�u��4vу��Dx��2�p�V�u�q\�;5�Nܦ�1&���[����~�z\��T�K��l�i��3�l�܉/r�E~�LX��z�' �3��^^x���V��BB��A��{fOvP#�`hK_H`����E�ڔ	��ֵ��˃V�(�ھ-�22�v�:^�G�aՎp>L�t���=DQ���.��ᢁJ��?�I\�hż��M��Ŵ$K�k�����Vm�#���uB���5���=�L`�����H��?uUφ�a��<�~��~���i��x�F��P�ơ(ZʡI�@ �<j��1�;ڦ/g�m�����e�3f��R*�����m�D��z�`kj6�
�ܝ�?�Ӓ�8m�<i(�������g:a��x�?�����o�j�{����=�3�`*OF�B��
�k��Ȓ\Ҡ�:�ǝ���^��%m/o�e��J�WM��汬X��Ox�\Q��\Ǜ7��֛N �A�yf��=Q��g_Z�L"��::�F�đk��I�;2����*���	m�LM�x�0j	�D�,u6��f�	Y+�?p=,ta)�D���,���z+�����I�tŢ����@~0�\�����!�w�#K̜��G̛��!;�_l�\�L�*����Ť�Ȝ�O�D�F��)�[xKhU�ȠSFD<��<�q����娂�s���0�#��;�� ��x�/`��E�`��~6�v}=�*�md��،@����l�_rK>g�y���D�E�C�κj�e�M(o��P�o���.��!�H�n�z`h����^�*�s��?h�;�1@>��zZ){��Ka�+_$� 5��,ycw��3 �XD��B]�y�E�f��&�]=�18����o9vrK���s��=�9^y�0�>DJ"9_�Y�1��e��d����:�6�]������Ow��~���K|1��4C�>Y�jC"ꕬ�&�'٦J�x�ӾXh��o��&L|�����s�����y�}A��~b�>*�U�M6�O�{�����oc]��!���ș�=0�%����j]_pU?<_}�4s��2�)��"��r�l�W�C��c��e1A怛���*E^#	�rgg)53O���
��S$ml�N�;�Ci5�'2ڹ#�j�is�f��:>�/g�Wvť���;�J�]O6�@�I9E|<`DI�d^�vk�q�~*���o�RAGsk~sY��FJ�{[�����`���i�99��VP��_�x:.����m��jL<��R�'ߡI�a�z��1�����rB��zL4����I��co�'e����U'��cIESڇ��������/|�1M�d&�"Ô:��pby�Ƃ}D�2m��X&�+�R�!�_�PḤI")�����&�4Rݟ�Uyk�|c��"�vr����b~���px�����6�s�[ٔ�a�G椯�����y]^?]�k9�=�LN���w&3�{�9�;,��f�eq���*/OB�w����
�<gQ��bq�z|�)��T�N\�$�Ϯ��:�no��Z��`c,��j���O�<�Ȳ�W����$V�3X�C�Gz�u�t�X��6d		*eo&rxC�s��~�	^j;{��*��|ڥ7x��ctЬuj�Hb)�davN�n. 6:��!b�{��iQ��bp�Y�!UrM�]�����50�j��=�K$�@2R�s
\��l�����]7.�r](�m �����&�ԝ�[�AD�ѭ�Ҹ �ve+���_q�br�m�(eQϣ�Zi�Z� �v���"?Q*�J�c�
)",),zq��C��䴢��eh��sPLp$=��#m ���77+� o�0j5i�-�g:X��T�2�z'�l�=�)�I'���ϳw��,��_N��:T|ox�|C�|�@톊���65��3Йڅ����"�����S]͘�A��fbUz��1)����W�N�|]2�S��D���޺&��w��ͻ��p��6�E���	U�D��!؄��z���0܅���qO�u6]��~�&"������*�F|F⽸�]��*��(S]�r�;�Ҧc�gS�X����JX�9��S�30���8�>-��V�{/g�e�5��(��滉Z/���iN�QQ�D(�{�������@����T��63�y�J]��j4b"�M-���-��?�"���+�ZƟ�]��g���� ��: �uJ��q�&',{������rg��BA��1}J]�i/ݓ����������4ܾ��,�}���+:@�.WMV�}��܁k���*{�ݝ��H\�3d��MnNE�?�~lբC�V�K�&m���~�EǱ�1V�1Yc���z޹��!k�E����l�GZ��%���t��*T�8�����#%�]�T�E�5��0/�@á���_|�g(56�����7�T�.��4���b��]��Ke���bៜ#�t?�$;�<�z5j�Gg:��P�Џ\۹j�u[�Z�sl��WG�iS~����
�7W;P5��i~h�&\�����R�FA�IT�D��vɓo2�i��o0�	2ñH�y@W�&��%$��d|@6��K�t~���Z����H��R�~�'1m+ZT���k�eϠ�U8�Z�6�ba��:�Xo�B�U������j�3�]l�"�]{ϝ��3�W�(������h|���HG;�:�ԗ��:��s�w5��OPv�"�1�Z:.(��7?$Ó$�NT����N�{_�5�1�����}|�e�)t��gK&� �^�:�{z�0�6����[r�6�"�ڱ���R˵^L�����G�t;B�Ih�<w2RuFb}w)�����y.=�1�Wjc��[~]�=84'3s��"��S^}̉i&�K8J6\���d|�)���H���L2g��5��Q��4B�?5Ý�B_<�z|<QŒy� �W{z5ȧ�S�`]?����fY�.�"��o=���]�|����m���cm�%=�R�c��Pgq3ұQ�4Ĥ�]͈�S7�>�+��Ra�f�ϱ3�v��DF;g�kĩ�>�fz��������p� #{.~��� ����`5��=t(�穨I\F��j97�_J=�.��������)�z��(l��C!˴�F܆;�������o��r��	d
ڤ>�R�L�{H��-_���o4̋`���*��x�3���ܘbx�2  %> ՘C�l�Ε�j�L�yF
�%w��X�r5282BԈ��2�N �ߢcf3S|&��x�j�զK�l�-�[�r(`��?�������~ ��¥�d{Z8�\.��Q��\b��8u�@���(n^� >�ǌ����M��fp��l=
���3v���l��= 
�*y��Edհ�v&���^�OL�?���D��b9�'b���i6�ab��~����K�h_|B�,[xg����@\��2�Nck9k���51��@�A*"�c�
�pm����I�х�e�x�'�j�ձ4.`k��+� '��Q
\���*s!)Ds���7�Mc�{K�^�\����*� Z��o�q�8�ev�*�ږW��{� ��#��F"�q��9#�A�Cm8�� >jᥫH:Ჰv�ܓf�M�ms�tE1���x#���^��\�Ff�aS:�KTV�*�q�#��{%8����)�c�y��o�5j*�P2�w�D�����j�fҝNt�̮%=�I��郄� *u�	?,���@T`��Y}�R�2��r,���u�K������f����Y]����%U}��������̘C��~��Ȧ��P�r
L���`��(�C`����9�I˸>`�yX�~�`�Y���̱����n9�r�j ]�3��L�c԰�0��)(*���w�,vr�Ǽ�@ �)��T��7IWD�0(�������y�`��SʵK��na�_��~%.�����%'�tR�n
��S�7�
�XD� �K���Q�(��t�vXؓkT`̏��Sr)vר���Dz�<��	�2˥�U#%��M@nK:�eS4���~�/0�5ڟ�?�7��'R��b�_�0�0D�E |�ʲ�@����c���K�3h���G��:�Pܱ�!��f��E5<9� Z�^50=�Y
�u(ʦ�

�8�`�e��ז$�}�+�p�#+�	o.�l`��)��tޠ��R!�C0K]f1͠5�����L��tޡ8 A��2֒�.�0Ze����[#D�}%QT�j�8�[����5D��1�e}�S��ϣd@����(�@ 	���$���ݨw#���,��i����*��'�a��p#���.��,5\�#�?|qN�����qA/�%@S2H��Qe!��I1��p��Q�L���f&���� QV����w�l��XS�ڮ ��,��GQj�Lj���R�{A�h�qS�����X�"玀H~Y��������=,��Ubș�o��M�x��Z|��/�CQ�J0�fH��p���5�M��:���[<�^�MT�@��&�;@U4X ����<�%x�!�Q��^���oG'�D���_å�}w�x�F�{�ţ�D~�kPĚ;�[ξ?q�M�̰Y������+# �}���U��h%���b藅Q���Љ���Qq
� �<�)]B� �q�9*�$#K��|*ñ@�a"gVǾ2J�詗Rh�։c��� N�vhj� 
�Ű�H&��-� J�f;�n_�^'��Ĳ}LJ�B�@7^b�rdLi��?@���ԀRЦ�2� ��P����U�c��sJ�9���C�=�&ST��<G�;��΄X�qRl���^���Ua&|U�e47�1�V�p�(���³6���gX� ��!Զ�������7�>��D��=����)�P�\-��s8E� $�����&�n�R�0tt:ȭ�,�*��Cb3Y<��� ?�0�(�GQK�������CO(#A��AJm�� )�2ՈA\�c��g���qg�};�0�
����Wa��;��9G�bOT�j�� ?���*C�x�:N��Qt�
9-�F��L� N!��D�w��2P�B)^}���Q�,�@�¹��F۵+�"��J�@�ܓ��X�	�(���BB k���0%C؁�QE"����cC�(�, ��D� �,������ƴx`���_S���D˶U� 5n1�c�Q0��w�$X�K�����9���E��0�wL�.;?WG@�7Y|�����]��K��g�5~�eK��	�e��q���������OD��s�y��=�&�@�Pz��$9I5HR�ZU4�����+�
P�e�YA�F��ܢQP��*-(��2�f�@	e�²�Z�ȴn�D����J!�0���l}�b��#�����q��˸x(dfx��<�ȼE�k���aڬ h�]
�0�VJR����c�!\u�#��ث��,�f	G�Do\	Lj0�����Z_1�S4-��]1Y�:�]�uPIy���w�vg�4�v|bN+�jP�UR��b�ہ�5#HŽ1�?QZKʂ��G�r�е�*[Pm8�x�c����v^%�s���X0� 3�-@�Ke!Ʉ�Y��FcEc9�ߨ��rK� ��A�)#�8?[��q�WPC��k Q�y��Kx�� �e$rw��ib
Mw��^���r�P��7�>��a�%^�U����1���.�*p�N�(��\@]W"�4E|b�b�׫�>�� $��x���E,��%h�
��յ��ï[-���V �ne�� 24����J!y��A��h�����wO��o�0g���p�}���&����3V�#l�����g�
^ }g�W?���H �1���ԕ�(���,�0���`\�p���F�v"aSJ7-�
i2IK���<����X��~OзK+��[�
8Łٌ�� 8	)�*��F������x�� �� @�  b\��(��"�7���3�B�9#�J&S�P��b5$[�c�j�3�j:G�-���d�_�R�W��B��T�f*�4F�3?(`{Ԯ#�����/��/���m��/E8[	v(�����t��MC��E��c�7r��:KlK���_[�Ŋ�#Z�֕ee`.pW�Ħ��H�p�r��u2]PDt�PUT1��G��l!���WI�Y��=��=�[u��Jmtt�����4⺰%R`���*���UNFV�!�<���S*A�rs�����P0��|c�DE�>5/A��+��w��DQ�'�` ^�hA�/��码� AN.B��@���¼Q*���Ǵ\� ��Uz���0��F��#U0��"SP=N=K�'�Z�۳?��b��^[b^"�q���n�^J��E�*ȣV������� ��[��P)�p�KE^S��BY@%1��D(2�h��A�`��a��G��m�K+Bb	�rz5�:��[]���~2��Nj:���?���BV-�
/b6�(�0�5D��J�r�(Ik*������P#�)�Vq%�&�b9���Qp����ҁvH���7�f�P�Ҹ����.Z��L>�X2�'��8���t|�1Ӭ��� %%W�����{G#��e��] �u�<� J��F���.�b�X���G�bpSp���� 9��RE�7
a����V������jɭ�O�Pe��a^����xZ�9,�  �A(/�� 4�P�,������h����� n5Lj\����P;��n�!�n*ַ�rs����:g���y��؜~qՁ�,x,>.F%+���|.9G ys���XꭹΈ�ߩ���Э8�e���x��@#�2���Ӱ��I�P�#��X�40@��g�r)�N�uʤЕ������wf�I��Bӛ�ԁ�E�8D��(GM�0,�� ()��@^� l(�2�NP�+۶"Dh�������qR(��i;��=���{���y�y��SJ��.j�T��2���8�8T�qT�.(X���ʃp8��"6=ϋ�.�I+C��J����@-��dwƬ��	C�sn���0��y�Q!o��SP�c�nH=��u%y5�W������|�����y!KAƻ��OE�Y[�6xzf�p<���d��`��k��� w������:Q)�P)���
������CT1}D���eJ1q�V�MP��� ��-�������v��*./1f�S��,t��F���h���}���MH�4��Y͹@|����]e�K�M�Z�aI�Fr\ݾ/=e'C��gr�{c*�r�<��Bf��>H����	�Y6;��ʡ��x�稿?�{�Ku:����߳�e���R�j���V-ޠ6Ep~ty�6'#���x����& P|�N�W'�|�2֏��ͭ������=�lv�_��b|X-��ed��"�XB���t�$9g14��J0�Sy���X�U������c����X��?���^>s�?��B "��b��1�y�`�$`[jT?l�(����m~�y�+V�Yx;� 4V��t�T�{��^���s��`�(�(����)��xE���^ȉh�D�U���;��
����)��")��*�@<���~��������BT�L�����JpVBv~����Qs�MҾߡ�8ص��ʔ�Y�PM���!&v]^��@� ���5�{��u������ �1��ɩ!5+�� �1U�uSM��=O?�^:�vz�㧼|���@�`��]�J�_�˭_�9��\c�eV�PEn32ět�u<��&�w�O�lf��o���h+��@�j�y!�k.�~?@�wC�����dyA.�R�I�2ͺBz���*�������x�l��\�����|M�O�F�����K�r�m��5�?�Rz��k��:g<T���48��DJu��߷]�Q�?kt�BC�n^=�����kd���Q�-�=K�qj��_���)��`$H$c�)�~�SPu�.�~w.\��A��Qoy������=o=~-��װ2�ƞ�]0�R��%
?�zW����6���YvM��qS��cꈚ���/j#0�O��I���h��?�>nѯ������;̫����'@������ Q�"�t��*��z~؋��00
��R��o	��;�[��c�Z
J�h��H�<?P#"��R�A�+i����R~��O������ ���ty�9t�7L�V��q+���A2�mX*nl䰡s@������ɚ\�4������%�r���n�%��^n1a;Jm�� ��q<�9�b��46�2��8`�ýˡ=��.%�IĶ#A*y�He��L��j�iAU���h�p7S�URud U�O-��S�s�3v*
��"���VR��.O��cm?1�?=!�c�E� dGrW�))�i�l������>�-�ߢ�f[�B��]��`����s1��q�`�5��D����gp�%P���8��E�4CR�E�`��K�*�S7/�!����7��w�TKJ{7�p�{��AA&��ظ�X��d�2������fΑ�i���bz'�f���.�@i^�ť�8����k�@ !�ne8�įJ~Lġ�a���3��	� G6$l�k�T���`��owN�����$)yy�n<��@��<ݍ��+;r���L���qs�n��m���#�w�b� �b@�$�"���rhB��֘��1��0��j�<��k�]�i��;x�I�R.�{�(���e_����$� ��	��,U}��?8�KҊ���zJq?�ݟ�@})�l��qp=�VK�5���@,{Fi
h� <���\�9B�$�}܀!x0����A���O����!������~,�����.,�x�_����2l1*ҍ�v�aPW�E���Ń�����@������.�?�d	��;G4�U¹[�^9�wb��%�	G(��`�������jX�1ȯ&Ra�ir?e����w�,g��%u��Kݨ�P�Ǭ���������)R�-fgL�A��x*T�R�˗�R�o[e��߉~%x�㦝��<S�~'�4�o�?�� ??�q9��?���� �hA��O�W�����'�+�M�K`�� x� � ���?�pl~4+��{�G� �G��PK   U^'Z�!�� �� /   images/a017e9db-93ae-45d1-af88-7a97bedfe2ef.png4�cp�mӆ7N6�=�Fnl۶m��fcnlO̍m۶���V}?��j~\��W�y}�� '�����o�%%D��}K}Na�A����k�sV�V=Ip���7IA�s]����ٔᱵ��ry(�A�8(("ۑF=�F"�*���$QF`��L�=���H�Pv�9e��sk���s�V7��WVV.O˵7\���+���I2�I`�Z݆��9����]��G��MXl�%�U�d��Yi����i�"�2�6`ZSfK%�@�V����;v��U`\C��;铺a
l���e����S4)IOޕ��[���C�D�����:�,?,n�S��j������d��0GOII������ ������w�����#;�X�"Ťh�m�s�=�$8��s�dؚD_3�d�??����TUW��Y۪�Q ���.�������D�QG��\K�h�xr��Cw�s�S��M�44���Ј|���f��\lj@�_�X���0ÿ_��~חk��F��ɉ	YF;����F9GGǋ��z��j��L�V����
��4�����������̏������3(�4�Lx�\�Ϗ�#�K�ۖ}�����}ӥ*�$&��ɉ+�����wMYYXRT�Tk�u�P��W,6�v�Gӷ%B�����W>��z��kՊ}���IO D��座����ZGGǽ�I�~#�&l_���4Tv"�L��]���@NW��.�_����� :T7�&t7�}�S�4Սo���J{��x�T�RdćX�9W�iQI	v���n�D&���|/���4��$D5ݖڳEb��`@��n��3ԩ����ݚ����u�ߑ0n#�wpU5~:
����1�n�`�χj~B~-������;� f����-�P]��r~P����oq*-��f���;�~ܣ(����(,.f6���N*4]�|����w9�޹x}8��>��,�Ξ�֏� J���H
K�Y�_����7x���}���4 �>4A�������C�qxuؿô�@L�K�"LJ��O��&���M��A���-IN,��c�&	�*��lk�:|�Nam4�1�#(�����ov5��wp�.�\d


	i�bP�i7Z�H^�6m���:�TU����j�$T����^�����lu�^t��iB�@e�'$��X��cq�A��b�o���!!)�9XU��a��{�|�^�3� �Q�<�����SWSF�￼���|D�
��ym�)!5^���=V������оA�416�st��(�	���
ÞI����x�X�u:��?��������@Y��O�6lm�]��z�MF�6P���;WQKk5�ю=<���8�-�%1�|>-�I�%6�;�FaDZ�t�{��h�L�E���E���2#�6����nLPE%��I6�n; �V@Mq߾��SW���>�xXO?ϯ�t`�zʎ \@,;�1c1_tֶ�*���������bF����>��<���5��А4*:zeK�~<y�܍;**
�w��@�8��h���v��b�h��y��I���rR�����I�͈�à7H����^<���ؘ����U^h�[���1�[0{��T�3!/}�b�Ԃ�=��<;:��ɡ�7�{:�еO�\I����QqQх�������7Y����g=]j�N�.(��߃P����-3v��yf,X+*+�:KKK����}��3rs��t8��JJI��"��ʂP�����B��MB�H���ܗw!a0<=�o"�s�I��:����KNnl|w8�u�X���2���!h��N9�v�O�r����h���l�ưQg<UTT4҈^��螮 4
�(X��'��c�T�4ic�c�k�8z"8j����ɡ�;�=����2�I�Ա&z

S+�S�}�
�QƋ5�Wɓ����F�gw�U�zֺ����<-����+�������qɴdH%5�A�Њn�C,B�����c.2�q�����r<�����h�6%�7��)yTک��w��ɿK�n���[ھ��?׽�.uKP��UHwJ�
E�)Z��:.Y�86��ԝ���ZHr���˭�w�t����t����W�?�2���'������JJ����}���yҖ���j������W�;�����������8����/��^Nr���FC� %�ѫ�\����Tw�*�-{Fz]V�UP�lLe��cM�v���r"�����0󲵵���8�"'��,�Qb����gI:U��Z�Ak�[����ţR�ғ����d"�w��"벑��V����[��k�×�����]fAAA�A�g�W��*6�ѓP�d�8X��ߞJʩeI���K�:���i�-OW����c�4���d����zV�852ZQ!b�mc>���A!c���� �s�2@3�Eh:q�x8[��U�+��P�~�TYY�L�\�~ �б�	����u}�5P/R����z��d��e��8Y&��0�g���u[�|HJ~]�;w�mv�yS�u�i�+�B:w�_2�/���춺>���"��|�w{]N�ơR϶-�i�15�̸�\�qEY_�tdj7[���m��e�۾�pe�����q@�\�s����Uk/W����{������H�e`e;��?d���>T�~��y	t�a�e�TDA�F;�����^���	�Y�ã#s��0��!,�-,	�}�v�E�Z��r�/M4�|6m�j���媍���,�����u�S9w2s.��	�	u��;�/��l���sz1�x�~����?|@��fMnJ�rR.�n��\�z���4y-9��D����`���MgB.I�,�݇C��joy���x�f~k�v��*������ә��g*�4���\?.~�n����RM��{���	��A�w�I�[��^k���q�����`�2���r�lOG��^Kq��SG�<��íQQny7�����F[3���~~���v�M�h2�~�ӟ���i�]���о_� �?E�f�)h-!����� ���Od�g�9oe�,�����⭢��g5@W~dr������F�CL��c��:>g7}�-&�e��	�'��b�L�$�Y���Z�6��Ml1��d����6W2;���P�0K�)L`�c?_���xw����Ӗ����Y�Nfr�DIӜ���F˹0:�.�G% �7�����5�Z�U6c��y�>;wY�}��f�������9uVj�,��nu��v��t������CB� E��G,����A�Z�_���'�{�t�f3��AKV]鿁.Dw� J�y>m���RS[>��]�F���غ�J-_�/Y�K�T����w�}A���x��/#C�Oj{Y1�m�k����߲;�D�!���w�.A��J�w���P�y�Gw����i��Zr�����;/n�}�.�_WK����n$WxX/t��,��$j&]�:���֚l۟;�3R�
��&PH �������W�l�k{�m�y]zؠJ���?{`"����<i^�ßi=V��hOx�A	�(��e?�nݭ$�_&�k�Q{�H�zl�p��ƽ{��?��={����Q�6Q���B�v�g��aZ���K$0�Q��ѤX�tʌץt��������Ce���j����q�>[$M|���t�rh~�n8����~��q���*S"�Ц2��q7��͠��Lr!P�[��.m�$@wB__�S\XX9���(��OC����I�2�ovx*?^n�%E�t�F��X%QU�9u��|�:yS��u�[��-�s��C[�6a�z1
b�f�����Q�:_��q[Z%���-��ا��5wOׁ���1�d�[�<6��6׳�6��h��������V�Mk���%����A�3F>d`,>�+��\{�����>u:�#I��D��ʩ��D���D^:���b�sd��<�S�l��Q �>^��L*�}WZ	*Y1�W���8Bn���Ukb��,g?��Z;�~���b*Brߎ-Uҳ,��,�}�?�͖k'%U��=�_�"�>qD2k�*��vAt[~���89,�C��c#{"�%ݢ�Xě^gU���O��rFKU�ڰ�p`��l^�ǭ���K	.}w���c<=zM��׸'�����X�yi1��'�pΒ�ez� G���9--�z�Q�Sp#ߡw%����U,O� /�Z��K�
^�q;:��n��+�����{i�1h\k���v�|�����;�!KF���f踉��L#�*����9_/�B��Y�x<�Hչ���'���m�3'u��ii�uM�	��h�Y*�m�1�Z���["�����#e�Q������!1���>������5?zl�l�Й�s�U6l^�4ق�q�7p��ΔT�v��i����dȯ�pw�G��(��K��v�r��
4��E��+~���SA�fS��9>���`<q�-h?֕��Ұ����|N�� �������NM��z�5��S��}�?ԫqD懿��S\��G��ä�2r��������"��OV\H�y�r�
~��ȷww���T�5C���ws�E   ��2���v� )��'l0���$��n��y��t�����oR���D�)w�䴢fӯ��|��￉��{�
��l�Ϻ1���鋖�Ti��AI$��&�����ɟ6�3\z�Irp��U��l���-�aEڃ'�Z�.�&����u�ݦ��ЖMUR���	*Vfk���d�f�V[*�	�PÌl�@d²|��dRR;��u?G������բ�v!y��B���P܇ƀ�1����K�m�pt"��E�����=�-�۝��$����h�u��@��b6�by��ҸV�C6��'��1:瑻�S����l�En��5'�wJV�'����q� 2s�i-���f/�"���[]M;'��l5G v��R�)��;����� ߡp�L���خ������3�m�Ws�O!
���������	��gȟ�V�|9+���T?�1vM Y+�r�.3HE+����a�Rz�IR9���#���^���k��(�J��kO{A��-`9���{�X�`w^��:-׻�l�x�� ���׆����~]��.�S�K�a�tp�?��SB����������P�Ѽ%�N~DH�#��ul۶��ה?��r>/�W��������BpJ��,�Σ�l�T|K������l�s���|_1,����*�.��U�A�ƥ������ʛ� �J!F�A�^�N]�q`:_8�K�A\�WD9���ct�����#\�48b��шԅ��c��r���7'�օ�VIk����漋-=�	ϭ���1$��o&���W�_n~�WTףe��R��%便ݦ �ϐ����=��j�j�>��e��^�G����kmV���7s����������2ؾ��TF{���Ҿ���}*�b��&��rle+�d�W�����b�v�-���u�箍��3�����V�ޓ@�'㔀����b��c#�rug�Jv���S�3��ph�h_=q�+���A�C��G��g���[�Qs���>/�g��湾�8�u	��ݠE0Q=a�H4L�+G<����{=e�͠�)��Jr�^*j���;v,Bx�u�vv=��F9����p2�u(�3��>�u۽nK=��oW��� �y����r��z\BudM�r� %p�9���DU��%b��:�$:5a�^��;��FdMY���:(D�E�6rL{xxxm���s*qR�LS���M�+���r��F���L�6��)Ir?�tfy� �fm��.��#rH�������k��j��r5�_BM��)v�lb����0�VK��(��EY;��1(P�AP�5�����Fy�����^[.g=�%���eX�X���=�=~�_���
�9�P)^e��O�g�?#s�������������,Ng���ɤ_R���B��:H0\9���T�{���r��!�� y�}~,]�1a��L�,Nj�x?�Kӑ��C�^�J���=��_H��6��\:���:��l-v ��&t^��/Z�o��D?��]����RJ.�<,,��u>���QV͡�Ǳ��Χ��6o/�KI�!H���"B�%��J���K�s<�U�w`���P~�Aˤ3[\��&{�&I��b�g����è�Ǖ�V�H��h��@����9��~��c?fݪ�x�t�����%���2��$~\�O��=U�m�:�����q=��O�(G���@�ח����o��Y� ˵��sl=����L��I,���I���8K7�J+���0��BW�vț�S�����ı��B�2��z���?}�k6&��ɰ���ښ��1�U&˚�@Љ�qZV]����J���a5|g��x���9�o]�TZ1iA���z
��4�~6Z��&-u�(<u^��V��5�.ڼM(���:�M�0��q<�!d{����m�/mg�6�T���/��%��n# �ᛖ.r$�w�:,�l8��iZ"�s6ۘ�$K����Irf�5��g�ʦ�������5���"!����=W��o�LQF@RX�&���	��a������_��U��Vt�ޏ�y���h��#�y�Ta_�o�K:β���.I�v�#���-g㜏&?���3P��y�Q�֚/�>��'9%A�-
剑_��?�I�_R�m/����r
�Ӑ�=����mP��� �x��C}K�f�1��PP�]kr{�x�2����or�1z�55�H&o�aRF4 y�ɚ�����+p��˽ن��:4�(���i�Znn�j���#h��Ҕ��M�נ�f�'��dcT�Gh�Nc;���+a8$7R�t���Y�����x���2�����D� �y���j��"\�K�IR��'�r�/D�XR9�Ujk�"}G�F̨�f��H�P�.�L���|��l?���d6�P}��xj-(Ԉv�33%��	2�#���C��n��eG�\�3���:\�`$���+ƏM R�v p�J{`` �K�^���h=�q����,� ��~��z�����,3eM:�Лm���pY�}�U�qS#����[�ˬ�f��5��%%%�8�Ɨ��$����rj?{��PN�J�/A�?[D9!�Yd-C����qs}Ź�I���(��[��әmO�r.#��;����VC�̛;�A�����p�-�ݻQ?d���D=,J�٤���byY`�,��[���n��zR��"�-��=��jkkV�Ұ�+}����h-�*T�t�4�� \��zx�ʡ`6\�@�O��_i7��f[��-�A�Á�R�o1�"��l�MW#��ϕ��'B��JQ�Õ64$�����{s�{)0+�N���D��>�'�<�s�(Uϋް��͆Ԁ�AV�}õ�<QB��^���$�=��l����v�;�zq \��#:ߙ���%;1�H�:���ߧ�Nj�\�B{F���w���[y��I�ʊ[	C�����7w �㡘����:݁�a"����,Qd�5[��T�{�:B{nȦ[�͓�J�3�l��+)�M�Oq���W��g_D �������~�݊N'��!x�o3���̱�GtFZ���u�����d��#eƓ��$%ݒ��46_��Qޠ�n�Y:>'��������Z�K��֝��U�3�6�aU�!c�.ܷ4���M��9u����6)���@9(�NR2BH��!��+h!���UX�~۾�VO�`�]bu�g�v��M'�T�6f��L	�C�ӿܝ���'߲4߻���긮z\�3]�����`(HU`j��i���gv��R�Ӹ�N�&�/���S>m�_����Ĵ�v���~M������囍Z��(��2Y�E��ؾc����$S��[W5:�{K"��lD�z�m���2�i-�,��K������=�զ���٦�Z$��Hs���r�yE��5mw�ݫ���[�e͓��RD�
#	(��}D�b��x����0���f���e4�9���ܛ.�f��\�� 
�����(@��g�w��m�/�ءZ�j�����'E�^��o;}��q�h��_ �Du�^ӱ?���h��:54j{�]_aQ�z�R��,���*=�����,���%�$���fTp"�{�
5p�<��S����������|V�V,�;� ���%��pbۯ��6�4|���"�PS�p�:n+�|��Ϟ����O��\<��k����s)�$��z~N.��k�B��|�|�U@�u8q�Q�={lQ~Bq�%5����b��\�{t��p�	�} ̠���"�J�R�/��`��,g��\��ȑ���I������Z���z�	)���BO��4R���6�n2���B<�c¯��*b��0�H���7��^�?�7�m��C	܋�9�'�%��ص�?p�q�fA��/����{K+�^!�aŚ�p�`������D1p�aW�	2|"�ͮ��4���2Kga�'Z����6�������v�v_�W����(j�Hl+��9֙~0���+� ��N��u�*(^��ڼ�z�a*"�7��@&HRC�y{9ս̔�T�o�#͵�t2�u��f���U'��`����$�T+2�R�����ŋ�;�γ���_A��+���i��Վ$�,ab԰�����9~ʲ�̟�'M�����>��'N�� � 4m�MЄ��j ��XYi�<�is2�KY�_ن��AQ�i����?�>�֝m�x�X[���f������Œ-�P�G������^�孡 ,
]D�K� =mk|QJ���,>�n�y:܈T>L�ڟ&/v���3ŕO�*��]�������^�	�
"���ף)	�%'Q��%��+T�ҷ!����)^m ?��܄��0�t�4�}�-����؜<�Gq�� ����א����7��[��b� C����p�*ܾ6pRZ5���lW����sZh�
��F��{�p[\1��A��J~}8�Oc��RQ�%��OH��w(��@R85�vl9���Z�'���gu�<LeS��n��B����i�ˈ�/v�p{^п�p�}��~��s�r�� �������?�����V:��3M�ɬ2�����ˀR�A��Q�BҶ��5��C#��tV��T=��`��,��&�/yt����#�>�c��De�P#ϨH�=���'����u]�!CbU·��\O1���	�դ�-Z�ݒ#-=�z�5�.o�jC�Y(y�N1����\_b^paR|�kI+pB��‼�����\�a´.$���D�ln��M��gF��C'
���Y�{�����ؒd�t}��)������B-���06�6\����7\��c:���v6O_�i�գ�^®{>m���}��0���7
&�y���˹���|@g�}l������Ґ����;JN� qc̅Q+�\ح�s�s��Ȅ�"��
Q�� i��s͍9�l�P9Λ�/a������t��j:l� �?{��Ж^uS��g�J ��;-��]eLԁPh,ny���-�لl��nےA�dxr�=�}�n����]=�v�*`���]���;و��گ<D�
7J+ta2	���l��Y��C���p�5LOX�A�B���2B�(.�#A" 
΋����`Ȏ̋�)��.��[F��*>��B�rbP��gz��ϝ��M9���^�L�	!e�HNg����
�HE*��vܝ|��U�4�e��A�\��$J�3F���ǰ���)�Q�*Qۆ�H��dS�Q".�2|�|������F)��M�����X�.�c��<
�o��1uKY�H�Q���R4T�M�r�
2�*�Q�k�O�7��$����3A�=� K�2L/�4�+�s���x����-���ˠWI?Vp멼Y��<�bڴ �L�6B���(`�t�dR!'��3tCH�i �$�ӂ,r`�#��`��`��CP� GX�I�/�ۺe�G�e��f��v	)��l�$����Ʉߴ�2�ϥ����)"� �Og4��#�bX�֕]��N���&q�ҔQ����v̈́Rkv�ƌ��B��q!53.fe������?�>�&��� �����Ɋ!���EQJ��5J���)�C�N#���@���}�2o�9I�,-��#:�`���(���B�QW-�����/��֓��O��^\L�q���Ԗ}c�2�(�(��ޞ��w��a�J��q�K��1����m&�E�,̀[���	'�[����zP�HW�����@|{{��SXXHB�A5��D"�a�?Fby*Ƒ���v��3��˝��c������M��Mh���I!,t��K->)���"!�R�&�޵򧽟#�����S��@�p}���� �&XP4��O� �4hޘŉSy=��ĵx������z~�#��:��#Ѧ���t�g��g�9((G��O{X�ÒL�v�3�"s:]ބ�������38�E��p"��Qd��T��]?�f��<�����N_v#~�0���qU)��c�D��1a$w�G� M�ӅHp�<x-�&�lu�{�m���)J�	`%���ub�ED���Ҡ]P�*���Z(���~��$��PeN�5��X�I�[��&a~1���?���\��f��7
/�O8wq�+��9��$�'��+!-k�Bk�1�F�0��pt<V����,�_�|!�#*�d艱n�I�?�d>�$���%�{" ZA
�|\�VqG������M�rV!cf�������O'���[>[.g��}	Y��&bI"լ16��Q���'�ͫq��o'��,|�w>XPO�x�� �]��{�R��Sm|�%$���$�3Ȑ�\�L:����G_���t%V�fn�#�;�0i�d3.ip����/�T�[_�aY\����������(t'���؟�ǌ)��O�`�2@���@�@ɋ$�0������%`��"�E��6��%��ɳx�M��t�Gq�I��=���WC���f�^��#z�/��w���M�d��篴F��3��P2�%t�v�@����m�E��#3��jDz�")�(D�aF:!��ʌ�V��r�D�,5x"����#�n����t�
3'�+T&���o�\�I�ع�mK�ǯ�������2_O�2�L�����UXqd��t��;\���P=6������y��oQD��1�4���b��,�/i00D���_��KO-��$(�y�Щ�陵��lp�0�A�Ĳ�kz���@��X�[A�x/�'b���}��@����G�l2/W�$ٷ����aD�,���d�+�|3M�פ��h�
&|C����:KPH��WP�����e�3C|���^J��r(�Q>bG"I�=�J�����=�(�X�����o]5�N���c� ��V�%���O@�¹l�]�c�#Ȓ��o	�œ�>�;�UK߉�����W������]M�>��P��,�D\Ta��F4��_�/�R;-_�xd�!���dLB���}�^�.��)��._�1җ/S���3㗒B�P �R�
����F[5���:����%UY�����莎��ӨT�����{(k�a��њ7D|����mi)8T�h��kj�D�;��0,��ST�"��]�6֟��)0���~"�!��N+�N�jJg��J⼜�1
I����ퟷ
�_�O[
�G�1�dn�t$tE���P�� �ez�V\�ېd��!i�,덅:�f�T����e2Q4z�tj�7|�X�r(�,�ڵE�fUin���M�`(�&{S(���h_;� �jz��o{q�������ҟV��� �D�2�Z�N:���O�oʽ��{�ސ��ܝ�_T1!j��3��~A�ܪ����2��y�&�6�V�Hz@�hv�G��41KEO̲.��A�^w��e{c����&��7E�Џ��H��Q�Z��눕Ԅ�v��9.���n��7?%���5=ܞnbc�a�Ҡd�-����Jԛ���U�T�KE�$��HJ��H�}f�"���怜噗�l	�m%��k��",dX�MH���n�$c�A�|L8��LeE�v�z�N��v��C�$�O<"/G��lL�m'��'/=h"�zڕ�f f{��Fp��}�s�~{��IC}<=2#�D�M����(%�iT�@��a_�j?�o���b��E�|5NcU��1-ʭ����h���8���:�[�V���m��e�I��7t�"���㹑Z��E��D�M=���w��`�#y�1�e����i���O2���
�ռy�$�8���z�:>⒬U�/���Й�3P�؈�׮�'&���Iě{����F�O�H��Ӥt�����	Jpۀ�whB��/ڠ;>���h�^�	Ra��%w"�����*�c�k��?c�����j�Y�VE��1"L���v�k����G
w�����8����`S�Π�&��B��4j�f���h��	~�Z��w�i�4TWd���p�� �wy�Y�n!����v=e=>)���bW����a�|x��2�W�����h1�A�~uo�m��"D���x��/0��V�z�KohX=�r뿬H�H�#3���k��z,U�ȵ\����9�*C���W2��B"�#/,|KH"�F�W:�3�N1��|�F}����ͦD��3]P[A�׭��s��3G����_J�e|��W����oF�|�ή��4�69""TFt92�$�)�"}��9��Q�H�k͢��^Ưg�x������nqr�N�|��Ϧ{D]T�O���<w��O��O#���CLF3.��K����:Y]{+�i�Ӏ��hP�u|3�;��nE�T�R��*����!�j��x����8��zW�}7�ʙL0-�����I�^z�0��]�_g��ʺ_��.�O�� �#B�%�;Cb6wH�vP����'n݁*���)*w��޿�+�k�.�L�E�X&��W����@P�Dm���ȱ�`�,����ؚ��a�]7�f���<ߗ��P���[K���;�;���(��oB��Q4����H*�xOz�����s�_8�s�P	����S�ro�{F��6�u��3���7bW���A�̝Q�k��D���E��柭���n �!c����F�\�b�tf�R��
���"LFͮ����
:�"z~a�����C+�J���6�y�����z﮷���$mh�i�:+ș�H��j��C�����p�^X��pL��bA�,iVm$�������)����7�������,�U�P�f�A���L�)��Hv(&D���f87� ��&&!y�i�_����%�����>@bzR�N�@`i�`"�"r�mZD��S�ȃ��游�62�������'���\�9	,��S$פE���Q{�c�j�;�L:�A�<v�6/oZ	<8��/��B��/jZwd�[�)���8q�nΟ��qkD]w����є�2�'���l%��ee��!�ftt������Ժc�ÅW������`� UW8e�C�����Af�(��b̴<(P0lQde�QV���0Lf�B�Հ���e���#U�@�+E��d;Q&l���XX:�i<+#격���)?BbTp��\X���H��LQ�1)z[X2lv˽h�ܾ�̕�8kʀ��������^m{>j�
���(V:`W�|�V.��S�1ӹ;�
��LSSS����������� �8�B���>s%Kn�a�+��E.3{�)�.!���ŀ��#�(-����W-v��΄7�@3���9�4	<�qum�!�:�@&��E�GGI����`tqBH�U_>ub�.��TG'_M4��ȣ����w��	�u�bQ3+ʨ�TQ���)���O�����_>ݓ�e���?o�6Τ��(�0d^2b4F&h<HE��c�{�R���r\;M@I����lΏ|��1c��O�4|nU�S1���֠i�S��F� �Dk|�73�ǳ��2�~Ns�%&޼Tj6LVW�n����}0����Z<�)����|�? �ϽR��R�z�������F$F�F��%����"��6����{���#����P�e�.�Q͏���|���#��E��hd"T&s��]X���w����+�OIN.5�D#I���^��v�<� ��M]��*i'�@����� :���}��K<^[Ÿ��pJ�fHMCHq���(�a����D��_�ׯk���W˕��lƗ���'���r�ן��D�x�r���t�_��A��r�����%r���d# 66We77���F�$�$�Ĩ�o|�K[I���{I�t�Ԡ=.��\̫`�pM�Lpl%��H��2r���3�ܧ+���X�8x��h@��B?�k�E��A��pR �ĝ%����wQ؎�>z,QO`������JX�R�:14E5/8���,#9:δ$Y�f5���E�!sK?���G��C���E��P�$�����Ph3��6����q� ֊ļ��S��3~]Cs��*[��F�:�����9�ϻ�87�T#!�� ]�u�(%��7��f,F���W���e�q=e�t���'�l~�3Z���Pu�S2��>Np�P��w��v��?G�1������.�����8��0�L���?���R��H$҂I�©ׁ^@ �C��o�vK�a��.W��	��#kxj�	ƎS�0 ��*�*�����_8?���E�`Ѩ9ԘW��p�	�&R�e�I�#��D@�c�BnG`p�Ҁ�S�/�p���Rq��8�s��߶^%`�律���t��|afO��K�)�	���d�����)�>C��9,���3������f'�̒�Ô��"�T�x\�� �MObI��5,z-Ü��w�y8�d�+{���Je�|F����`/Dx��f��L��(�����O^k��s� ;)V0�v�^+�(��W,������bB-��"�D������ay��.da����CVE��Z*�h�߆}���x��L�ͨ��B̬��� ��!E���@/8�|}6
Rg����7�:���>@�Zx)�&���<�i�������8���D�m��m��u9����2�D���{~8�-�`}�w3q�$�^;h���?����$)���V*6��.
�(��M�6�G�No<��:Z$Su(N<���O*�^������ݱj{�+#�+G�b�����j��8g�����3��%���"GUz�&��hk#
�V$@Tp��WjK�������GOk�	#eA�;�@��E��-V����ah�"�5Z�9'8����C��`�?W �Į��6��I�"����k�g���d	y��j=d\�'W��e8�`VK�șcfǡ-_MF�>�b�#BF#l1��(��A���ɮJ4S�=�Qi D<7��ք`��%;9;1�d�I�L�cU�U<n���(ߖ�6fp�j�ur��i�P���|Ս�[RR�_h&ǢZ�'l)H���p�����X 0>Z`z>�9`f~�E9���v-�[L6o����N���䰚Ƚ�� ��L��C?�:�K�c/�-�rk.x;�p�YԴv�&%�3��e��oLu�7�������� Ǜ�������v�o�.ſb�44�����˘�'~r����y��II�X*�aׁ�?ow�&���l�Z-\6�����Zb2�	���m��Nd�n���Yu|���ٳ�M�ɔ�10Pb�Ӳ� �_6ld�z���\��XSN'Ĭ�h������Pm�� ��a}<U\\KUQ��̄��
�i�ٮO���9���������	���7����9T��*'w�����n��返�ޛ�R�9��h��3����*����J�ۅ Zq9Cb�`��%�V����饨�@q�|�)�+��{�+bn(`D5 9��Ĥw#Fw?�/�d�Կ���X��k�c���y�&�h��g-E�.K���٩E�}�]�^i<��$a!6��.";S�V+�FqHd��VM���4A�#��]�2c���!W3	�;pv顽����t%�+�(�
I��h-er�'J���4����� ��~�D�:t�AQm�1�{�2h53����SW��o��ݙ���h��=�7�]����>�_�����i����{�E�P?0QeM\���!���g�?�7�x0�vIJ���CR��B��	��ԆfU�Ԕ+paB]�E�����	�$�b��5.�uY`��I7H��at_̙I�K�O� ����;=��a�tQQ�4�܏����I��,�<���.S�l������kc�^Oݛ�C���	�PXz��c���>�^)�ү�)߹���f�\ķ����19�oy,���k�e�E�� �D&{������Xtӯ���BH,:g=�9@ƿ{��M.�\��s"B&�W|q�����,�e�=�~Zو_�ȗ��ݓ���U�Vٱ���!�<������`�n�Tәv���R�C��c3&�#��k�0%6�:dj�aV�P�*���FT���kMO��y�B�H��RH.����S���X�-y�A6��:b̖�V������R����ԭ��}9�QZRIQ'�6�)�ڵ+UOj%5�
�[=�/!�U�<l���^����`�ԣdS��E����/�Ĳ�
�׹Cm&��*t-e��0��z���gOV5�"��]�4#�A����,EN�&��W�y�J�X W�6fΜyzvv�ffW-O��S����|����J�[Ǳ#�2��j}���,�PRآ(��-�9���:lp���ԑ��ssSGaVVV��v��sS�,Z���/��F��e����A�h���u݅��w#�FB�B�(�M%DSfA�Q)�(bdbh12�$�J 1�(,�㗲,��4����r6�)����U�v�Q �,�b���G��!�
~۽��O��P;#��Oaq)+=l�I���������Hί�m{¶�:Q��Ea*�p8�To���.���!S��##�G�o|�H
2"epe�w�S�֨Q��-4��3�<t`���tŗ��AR� a�� �7Nm��ǆ	6�9���3g�9����^h�$b�S�΢�3g��>�=9#I��]�Y�{�.�Cd�=
�P�sоe�¡w��U��h�̭I��n/���*�@q�����ؚ/�<��l��J�Q�05���0��Y*���S� �A}�k��Ʃ��Rԓ�M�!�SQ*�C�̣��kC���}�\�`�B�Kt��&��@��Տ�g}��)C�cC}(��e��/))��)oii)�����'� Ŝ�F&�I~�A#d�q#
�)6a������]o{o��r>e�Mc��v�-�T�}�Aa$#v����X�	�p\��~�wҨΝ��=�����DD��LEI�`��?A��R�kZ�"�c�
_7an�.y�]������kp�ƍ'����	����q�B&�+>���qoe�)i�s�e�!�aHj��"��t�/t�z�\�$��j4R��Jp�i*��p�=����9���7=�ɏ���H��RMd�	��hB"2P#�r�$)(++���ݘ6�|�~][�;�؊ �� ��6ΤSb�a�|�n�ah^�"eC7$���}��(����o�2{#"��#.�ʡd�u9��۷�p��Ә�<�TMG��:ؿ?�t�d����[�) �$��<\��K^��#��Ü8j�)��h@�I��%;��&�v{y���G
z�d9�0Ba�?I�����D�ՊM�b��B�B8���/{u��G3�ϼ~�ʏ�/�NH�d�@!v�8��?�F �V�v��LX>v�U�h�����KCV}��8�J�<=�E��
N9��G���w��uLCH��0�LI���"�C�R���5�K���ڮM���O?uY��N��u�rdC�J���N����	K�7|�ë[�џ�(�e���$�v�*�"C9˷��k�YQ�,��+N�?�-긶�CSNu/��0�hD�SJ�nF��2$[���jT�.:PQPb�a�~	�gވ	?��7��ˤ��X�H'�����%��}��d"0�;Sw�233��������E��MR?��HegS$�L��tjw݂g�sL3}�E���;*:꒓�K�r�8V�	8F�cR'�H��p}���4v����6=#@��n��6|ոG��S}GL��o���Sp8��fe�X9b���P*�I&6=��M�N\6�qkz���f���ݸ�����I�	�	-�{G��F5�	NBɄ�LQ5E(�D��[<DnY@�h?|N~�^�K��m]7}%eBaqe���%BDb����߄���7%&��BTC.I����.h�^]�](ڽ	zpe��rKPe�բ���Șo8QX" �X~��$�?�|�f�܂�QLr,
<h�a#�/��Cb�
���$��N�L� ]m4Frr2��ˊ���B�C�C�d6>��Kv*�E#�h.���<\����?|�[��d^v���Ky��J,�|L�.�H�e�9#0s�;*�Lf\6LqO65b�.��9�����N����II_˂)7?��߾�4�ˏ�����p!� ��섡�K�Y��0D&!�Ѭ���ǎ��x𳮭z<�⋯�����p�JsUq�W6l،�7���ㄐ�앟�yp��9!�����<wD�H���%�p�F8 ӈ� >I4��n`�D�-&mI T�,f�Ij
�}�PL2�Hh2�&Bl���6xl@�	j� +4�FK`�(�ۃzi^xm
c��i@�p�{{Sk12�W�*{Q4�:(��H$I�Cb$@I�A$��x�g�.���#%%L�EGZZ{��TrssQ�Ĳ�J�n�$��O�d"�0/0��x�v���F�SL�t�ێ�Q��[ͦ,\�հ�m���~Z,Q���c����b��D,��1Y%v0-#������ڐb���
:��]�G���@#b{�w��Bb�!K����͠bf:$A�B�^��D�*���D&u__>��*I&�-z>����z��빚��v�}��#
n�
D�vH2!��� jZ�'	R�)��a>Q�H�u�/�B!LQ�4�'�b�(��ah>A��E1v��Hņ�����c3� Ų(�Q-ʮ5M��/I�C�z$I ��~i\���I��ͮ��:y��k�f	�# >AD�$IB4e��6c��g��7�$I���jnA
Q0u��XH�ihA~�D����;�9p�@U��{y�Iff�����������Drii ��X� ]u	�D�X��i�e� I���؋y��(v��E	�$�j�+�r�i��i�~QD)�G3|�,��)�N��X4M�Gزw�0|����A�9��`0h��7����B��n�����~��&M������M� ��n�I�ʨ/��,�lARu�#�b�դ�@�(����^Y����^A0�h>M��J���i��;~�gw��dC���cdBu�)-�,۬�Ն'	�2ʺ��t5C�����A�C�NV� ��B6Ð�(S߇i!Ț2�2E�
]�R�61�P"p8e�v�<�(��M� P,�TtM`�m�b�&* �iH�jd����0o'�z���BWl�S[9��OI$D �>�����!&���f�޽�vB^yE�(�P-����9P�w�����S !Is��A-�Q����A3G�=�p���io5^��'�~�u�B��6dW2J�.AQb��!��Fy<f<��s+�Lt�Ȕ�Y��J#�nR=}Q0��ӡ��n�x�A�@����4U�*fR>1J�B+E���6(D&�ę��NZ>�;�Ye���)S���$����Jb�yM��\�Ϭ�y�&�I�����`�2p�,��+}��⯭����-�|���׀g�G\&k���v��0�w���H|h3�O��9��{�^�	Jc��J]7_aa![O�|"Lڸ�k�s������pJMM��I�"_�7W}�w��C��A���4�d�P;+K�b���v�2e�աkad��t����XZ^]�E�^�C4��
B:%nT�zK0쐨j;�d��Ǽ�Ȯ�v��۠G���� ��,����Nͤ�� =�RD�W���z���("%@(""(RC �^�zUT��`EZH�����}v���~{Ϝ&��$s�'�L洽���w�e��-#4|��b�0���Dh�2��an$�x�^I��t�"�fN����W�ʓ�E,N.&���sc�^�W&�����kxLӧO�M��W�\,��E�Rr�AU�N��~�R?Ҧ��c��Ӊ����&�L���~��M�OJ_���Cִ������_i�+L�4���Σ�q~
#)�t�[�w��v��)�$R���	�L����_���tI���H͉' �>Q׏7�_e*2�cQ��G5�#R�����:L�Oq=聆4g�{d�1u�Ȥ��LNu`�p��k����[��i�$]l�=I5�;���$�� N����#1@�}B�`�k>0�6��ocS`�f>�׋?@$P�0'͋	����5M����j��G�Z��`2|}�5���Sʴxr<�|}���7<O�$�$疔���O j���[Ln���/�|��7121B�X�����ٔ�@bC$u��D����4'����f`�p,l�� U��E[��2b �Ж��X���*��aл�ߘ.�8o���a�XQ�H���>H�@7a�L_�i����Ш\������Cխ�gd�9ٜ��+WxdqPxq]?�s��?�����U�K7��-��ZO��q�8���5lnx�la���Җ��ZE�"��|h��L�� @U��Bؖ# ��Յ,�Ι�	i9a�')��&
�����`Pp3�_U�3���}����tL�+O�u4�g�t)#N�B5���Q�#�ۅq�.�F%�,Z�����3�Hi��@0UG%��>��Lb,k���Ņ��$2��=��o��?�>?� 
����'�@��q��C˒�u�5y#�'���?�.:~�#6��'�Glm�m+�N:�|�MFoGʦ��ָ���N�8q��IW�)�I�K�e�8cMy�q~��G���L�Ɔ�RT��ih�w�����gd��	�0��
3�oC��+E����g�(�\d[�5��*"SG�� v �UX�)y|/,"ې��>X; 6tv��dRr��6�9��/�R)����R\x�� Se�$�
	:I���l.�R�!Z�'��f��P��Y�{�3B#��|Āʳ�8#ߛH��AUH���ER���&V���� %���L�-��8?�)/�$�WѢ��/���H"��jmU�b�ݲC�R�d*�t ���]��
l��쉋s��c^k4���w�7��z����R�:,��\I���ڔ��1&����I�o��O �6}����#�K�D%4މ��ؾ����$�%m	�"�HE(ն��f$�!����o���z�`�����r�N��u���{���)W������ɔS�ru�ˆ|I��w� ٌ��i� i�q�La�������8j�!S�L�ʶ:��O���4"ھ#ޫ���$�3�z�J���Xz������]�`k���j��\�A}sv:�5k֠�SDSCl�RB_r���ڵk��A����]i�t&'��ke�<=C�a�j�+��=#�plS���Y'[�����
�ȇ�N�g1]��V2�'������U��i��3����6��$?%��I��R)�7.�%�gυ��dKSjS��^u֋�f�"tj����3l!q������IIH�9��:���;�ǜ]&.����&^}^kk�9�f4(Lo�_��K�#���L$�R
�Q{HelF�q]�b�w�f�Ү���J��:u�QS�Q��ښLb�_ke�����I*N��ժ���D���y�k"I�$9�Drx�:~S�eH�������Z�ʒ8��Cf�ױR��J�k�Н�G�IJn�4$}F�Bg��
"tژ�S�� i�{*�~�7���6u����ӷ�̽��(�H_R� �"H�T��z��0D�j��W�y-^�0��Wr@ ̠�nl���w(�k���o�?s�"�!.&Sq)���D���#YYN*��r��E��Y�es��K"-ύ6m�tٔGj���Sw�31��?�?�����2&���D�v���a4+�C�����燼~H��:s���n��zm��y/����du�1�lXS�l��%�+!�IZ�� N����4�*�5�	K�b��_��n�w-Z��ܶ���0��4����9�:E�dl�<��-�r��T�ǥ��h�'�a��)�j��H�m����_�nU��7o��D��M?�z1�]
�"���#��Wռ$�jVwu�E�9��[�4<�1�)�Q(U�U��tb鴑eɴ�$H�Q)d֭��Ea�8�[-������n��bf$MA�HX���1�C�_Ϧ�X��
�C���\x�X�	ؗ`�K�2xՠWC�-[����FD)[XV�E[K�?��;�klo��K�H sP^�g	v����~I�-�ы�MA|	`Lv����+�jZ��^�%�̟����{	���"�oU>�14��>�Z �+�9�E>ecRK�D�v�C5��!啎�^�dI�V�Ā�-�Y�I#���)�m��o��o�/5]�H��_ˌK����,���U��Ѣ��H1iJ��1#A��Ŋ�u����+� 9�)Tx�u�DI�W*F�8p�.�v0�.�\w�c_:㲛o`��*`�=Ҵ��BU��V\��k�E���nFhhj �&ʮ���^�%����^��IhM�I藃赳�ހ���}ī��v����+�=�b�5�Okko�o^���ݱ�������J����L�4C'���
R���[[荒��t��K�3�KX|��X��6��5Y?:[C�3�V�����d�(~$0aJ>�O�$�I�Ew���5>��"�Ӧ#}g�zfs�l�Œ�#�l��٭\׊��Bӆ��5d,��F�e2���!�x����0	��"��,"Iy�*GH�n����=�М�I���u+%�7�U?Ć=(�\47�Hx�fWO��傛Z��W�=��뻅��j�d���_{ϕ�����o��,�f�I���
�0uB�i�Z�\D.� c��=m�dL^���m��bjD�P�U5�E���t�ւ��=�i���Nr�;���k?���`_a
;R�>�mHu����e����`M��y2��`ѝm	����e1�y�W�[��7�>����p�@�� �qڍ4��](����vJ"���������Z�k�}�}yޥ7߰m"�Wg��w��+p���㘓Ne3h�ס����Ĥ�T�Z[�AO٘0y��R�G� �l��a�"S
P�}��jm���2L����j0�e�u�\1��Ѷ�-�����+!_�U8n	Y�D>�¬iSD�aǦ��eƍ�f_�[X+c!>�SKƢ����h#�E�{T�R�ю�S�:?��l�zdRi��0Vd�$�^3<�uYx7���%{"�W�P�zŴ�td�0�6��	J�GWv���+
v��a��`e['6�Q	5h�#�FƤ�3�U��֋LF��A�C��Ƽr��/�m�4��CO?J�2�9��o���)��H��6y'�i�ꑡRJdҁ�zH9��3�(��C���(�Ͱ����Ղɜ]'�p��s��V:�-9��~c]{ەI
�Z	V��q{1���v�,wJ�=9��)��\2�SQ]U]U��B�\��nm�2�q��k��o�Y��_3��?����N�\�"E�&��A��'?�S�z�2`�uS��k�@��~F2�5����S,7�Ѷ��Ӌb5��EZjMg7ڻ�P����Y�t/�%V�����m9�a@J�0.W�b_�\P�r�fhj'~,�+E4�4��ԏ0p�D�r�GɕsR\I]��]�QD�e����H^�u�^`�ma~��7�s��[m�sV������ڶ�rz��"5��+��Oa��z8t�_�['�of*J�JJ'f w�y
��+�oT��ǰ��t̀��Nz|��i�"T�Ҙ�Y#s����E��"tH-�@&��I6�r���    IDAT��Z��T�F�T��H��5 &�p�*�k���PI]q?�T�Tf����0�u�,����}e�$R�i�eQ��&c`7�ы �^v�:	(���+�F�Z&��kն�Ux޼�M����!��Zș'&B�Ag��@�t&3�b�K��7i��!��Sl�98
n�my��62��	7�s��/o�c~-߽`Ѣ��u�_J�!�J(���]��,nQjs)�D>���-ӫ�oR@3�;`/WR+Yh֊��J?zh�1R뵜������6<JcD��k�������_P� ��Ȟ��;���c�b��0��z�F�N?C_#I����>��뢻X�zJ`��v���}U�j���2���i�Ismz{&r����Fv��U��r"v�T���+�y�Y@�����c�j�t|5
э4�;�a~2^Z݆�~x*�#S�C����IR��H����6K/����Z痊�1S̓�%H��I�<W����`V9�S���e���^qڗFے^�h���?��_*
�p���ڒ���!�.�S���T-�6g>��H�s���f��F,�����D(b$wpg(Y���9��cg1��\f�&�H���^�\#��fx������*ĉh%?��'u��ٵ6�Z���݃r��L�h����|;�BU�t>��;�$zX�"&,Q58{���\r�7�Ϥ�ޗ��_ˑ�����0�*t�b�2T�l�a��KkD���[7O��'�;Ej��Y�N�����妋���Bx��<7ڬ�V:��_8	�|P�M5�%隑�LF+�\�d٩mm�~h�4����̖FL�[��!���(o�x�2�"8���s��M�t^ǎVb�"�X7M]�����#ӂ����'W��iD�$T�d{*��4��R�o��5�c-���f�k�LޟL�L�U�>V����^]k��]�+��4m}E���:�zJRbL�򱝰�6�ܼAjujX�J�@�8N%LkN��������ѷ��p�����8����&�%44����~��]��0���5�Y��~��y�c0Q�Lj���]�^��!�.��n4��wh�$񸶗�䪥��]ߺ�"
�X�
��7`��&8a���'�}.}�Hl,ҫ��a���+܏�W���!)�D�J�e��g��������k���lT2��4_ʒp�y,0�JedEkOj#������"�$rJ��D�2�8���V�~
�������S(��(���_Z�7Ry��HI�(`�\����+�� Y��z?�{�����"zW=#:NZTB)�/6y�>粐DiD(�h�������W���]��Q�Rh�"�"���4�v!�L����nj��$Ə�+A�a�;��v�����e��\�n�N�#��}�xLn�����ϥ��f���C%??r�u�� ��~�XC�c-P��{̍o��$�v<j0SW��,�$*I����d�Y�Xg�P�$��Pu<���o0��[�y�?��v�%wM"hYT�:c�IN�XSS�H�(z$d���~ ]��j���~DV���ӷ�D&�+�An0���Ⱃ�&s��B�ђp͹��mM��*���_�Ҋ��*BJ�����:��%P��e�����3��˭8���Q4�P5�pC�t�+-2�0�������	��D6�Ԥ���I�VQNe��Z�����W�/)--��SwB�c��}�Ҷ#�uh�cQ����(U�P�����t��.� )-DsB�H����cGnZ��M�\S�'LkY��GJ�Kbw�ٗ��Ex��Y˥<I8 �8��qh�Jm�J]�M�&��K�'c	)Qg��C���A0a��������y��)���(Q��t�$���7�~�`Bd��[��Ɣ ���"��V�Ѭ�����RȖ���'� #���oR��14:�4Gި�Bv9h���܎o�����f�����|�	
_�d���Y~Q�e�;�l����fx�dc)��l.E�T�^;J����`r����]��<U�������	=4֧d�g��Yӣ1���5�=%bD8ѓ{����0Q�K)t+U��>��lN�&�Y�x=d܃R�#K��^	*��d
��u���+�en����D��ɒ��L$%2UK�W�u�EA�ry���M���- �]���V���w��w��d���4c�Τ�n؀�_�NÜi����X���P�]�"ϴ�48lcj���53�z��Q��ᙕ8��K�^�������I�TIf{��^d�1G-����8��g�|e�������l#.��b%�ن=ȞS,��i��J�fْ�]���C=��0*�o���R)�d-�!�Hc�#�cK�҇G(�
̀�qbW�&�Pl�)�^��\����$�.��fOj$�=��c*����Y)�o��)�x�����U�^�엾�$�$=_3�� �{�dE0� Ydm����>��
ձ���,z�� `R�#i��fR�̯��UЖ��Zv�S����E�w�Z�c���Zg���ױ�B'4����EpT�����X��2��'�O7���p�w��gP�c�LՓY���� ��i[,Ɠ�����6����%$@�m2�$���+;f!���iźR�Mx,vJ?�Y|+��y�A�L"�ё��0g�	7�}���3Y�t�y�[W�î�:���w�z�M�I�&�<�S'e`���+!G�$�7;F9�>f]а��o¸�	0���FI	oj���h�}o�q�0����1�/�iC���l������6R�c4�ݐ��°/�=�zpc�,�k�D/Ӏ�сu/?���KY�\������:Dكvk}W��*�]��ɢ�U�c��."���ɔ�������0�yAF"����s�U����с3f�lq���*(�v�65�UJ�)�Q�1���KR��Jdmq#��t0R���}fO����棯��M-x��'�����\��:&����=ߐ���]�S��u��4NX�{����ݙϤL-���a���_�y׊���%-��Z�p�f{�Y��m����)3�R?�V��qQ�W���O���u����aVK�3���__u���3Y�p�y����Da�v�w̘��_ASC�Mc��b�Rz��\9��i�����85�B��_�Q��53���<X�Z "Ug�\��h�o�|��Վ�s��3q�_�Z�+�6$����N�0��BQC��6����ܓ�Ψ�
�7%����Q%���|�El��g^^�^*}�)ɬlU0���ǿr��7]�f=&9I��A�]g^��Lt1#�;�	�Z��K/���@5�ꡧ�_r���s__A��e��=$K;l���w2K�9���%ؑ�#?�^�z̿����ܛo�W��n�"Nv��8�w3E�-ޟ��j�˔�����������%��}⼟����˵,6sR�0i8�#����l+~~�+�w�W���?�l������L/\z^[[�9ATA����
J"�8LT�O�	kHܣt��%O��Dz�iV�
���)�FL�� �pP)�H��C����"�$uyC��=��
��۱�$q�xeUT/@BG#�PәVGA�Z<���Pg0��c�*nL���Sbx����G���+��L�ƙ������W�]v�uo���";���^@d�����f�A������%rhmm��fΜ)��um���d5�.��L�塏�`;hD|�<����Y�׏�&g��.��5B	/)����xbm~�^.��ovX ����Nͭ�B�VA���������M�V��SO�z�u��?���]n=�B��z08��ԏ:�Ҷ�ޫ'����E�?���=����dF��w_}ƨ�L�\�컭�mg�&2 )�*B )#���>���0Q�tT��;:�Zv��x`52z��{�԰v��l#I.���]�^c�0H�$c��,��}tvv��A��-����cc4B bX�ב�͈����PC5�F�%Mzj3�7���9t>�8RZ�rQ�4N}�I{�s�,{i��6ݲ[��uU�>�ۏf����^���)u��������N����ʪ,�{��ԑ��I9,���s������oz⥶/R��`r��q7ݽ��Q��52�TTdB������IQ��A�EҪB����*��=�; hjQ^��.�b�*�~U�A��B86b;�3���-���>2���'�<����ڑ	���v�|�l�=][d�]�|Ȉa	r�Z;�%J�q>_/j�|��rL%���0�nd
=k����w�}� k��:�ǚ.�^�EJ�������Aɬ�=�!��[����W�%ZE�l�ۏlԏ��F�-!8��}Z��w���r�2�4*�>��,��0�9�����`�.���ھZ)��
ڥ����oo`2�$͊Leqm�^�,g��h���Q��Y����a54vZ����l���dh�D��7OM�^��[�<�{0��'�:����`yf͞�
�&�����u*�D��������,3�W�Z%�x}}j~�����7��+���+6�0�Ër����_X�䟐�հ"׏��iW�g�'����s�ߊ��8&<Nos�4�ȅVlC��F��	7ȨY�y&����*���ҡ"�۲���cf���S?��Ï������G_h�#��;vw�o�}�^{~[[�YC�\Id2L�,"SHDj٨Ɉ3��^ �&�q�����`��ݧDj0��C\x��$j���c[��v&��y��]~��7L���I%e1����
h�v��Ӈ�ӧ���/�M�`�<y�D+]]]��㳞A�)*�H$Z\��(C=�D,��F�����l ��2V>�gd�~�+����v�5u��,<P��*����ܖo�w��)tɇF��!�V=�{�J�
�Ђnv�=> }��r}8�!��E���o�eL�3~��K~�Ly�U��|�ع��_�?��7�l_�7nL`�㣆�t{�H���4D�	��*0�d�0i�,8��$��3���a;�4+Z2!4�r�%J�$��q�wL^�u}������7O�6�����`BI�4P)0{�l�}���M:;�$J���Q�\�n�D/���"q�t�#^�: ������e"ݰ����C��7r�R��;\+~�TT������/HG�`r;�*`Rv�L�7Ay�uV]�%�����h�x�w!���v����OoD~���Jz�D�4�� (���=�L�F˟��W������G^h�
����w�w�揾�[&l�e �X|�
Ӧ��b�!�0-�f�h��)�����S5���W@�v{m�S����10y�p��޿݃ɒ_?9���7��0aAp���d��}Ҁ�A��*����"�pƵW.��i�mmÔ)S���I�I]�,+�����gv�����ZÆ�n���U��X?��ה���'�<�g�~9�@��~�n����r�5� ��x�z��k7��[+於f8 �*���%�����Qi��󷶋}(�z�LU�"��TdȆN#����X����3K����Л�K�IF��r1V0%����;.9d�Z��W,{���G����c���%�������[����EK����>oci�D���˔k&�衮�����jԍô�t�{���PȐ���:��!�10y��ƿq����{l�Y?���-i��#)�i�h�f�o:V����֑�U�؀��R�0i�D(�W��h��+F����#� �⪭������>�>#ޔnh r��t����p�ͰP2rhG3�z��i��Ŧ�Ƽ�u�1'`3��U��N}5�W����g�0����p|ef9U�D>c!*v�^w1�,Cw{`:Jfϻ�B\�e���
�
��XPfQ���9�����W�L�u�e7>�r��X�J�������y����{�=?���E����8�4���#�A0�L��q�~�a��(0�<���O@�D%
D��d}�"�m�S�{0y5�	E�F��ׄ�R���p������^����"Ȱ���C��I�ɸq����/yu2��0��:���W�y1�v�\blO����n&�j���*�z��y��8���� �,%	�7�/�����|7A�2�Mv��6�>6�p8�Ԯgl���<��9p�2��c�}C%&�qR�*��"�f���>�}2t?�e��,���q���&̸�� i*�����"r�����ڵ�}������{���)�2���_/�w��5��۷L�f�⻀�
�#�L�c���#�T�ʺ�0�/�I���c`����x��(R*�ʑ<^Q��'�1���m Is��E�;ڙ��Rv��/�R�!�.��T�J��Rñ8ˁ�#�Qj��Z#,�V͝$��aN�}&��&,-S�ηM���w�r?=�Ne���O྇���u��qzemQ���c����$jH�0�o�M�_�kk�?Rjmxʬ(6�$� )BS�#�b�[��_�vjɃ���jz�7��o���O�.mI7��&�*��s��ѽ/���Ok��q��cŦ�o�{�C���L�L�E�7�q���}�ָ���g.�f���mg֦��A	M���+�9{�d(V<'^J l��H�����\	�p�r_+����Jm����4���Y�}��V`��~��Nst�-Is)m*�������	�=� �0�\�lF�#�͈w˟|}oo� ���T���i���?R=@&��R�1���W�� �aZ:�rF:#�0�Q(�+ �I	9�I��6�l䄹�y%d�)x���������d�`3��1�������j���j��W���ּ��f(@4�����'�x�x�Z���֡;����Qok�`�Yb<�k�EU��2l�GX�腅�bh���"3��\��ǜYM�Zp�v&����.M�҉���a ��� ����^���]��L��f/P�����cK�7�5�=���4���X1s���h�)�X����"c�E�\6��q0,+V��Z
k%Ӧ���5k�$��H1�L�0�HRg��bPc0I���Ӛ��@���B(��X�v�r�V!�WE���ǈ�Qe+<�N�H��D��́�p#���4��� ��$�>Y���%�W�ު���dn�{���椘/�k���:�(^�w%��M��j��b	�tJ�'mi�*E�Yg���A��5��҃�Ԭ��W)
H�Ȱ�@ ;+jά�X�+`r�얫y�Y�.͵��D�	�ʠ(=9�UW��G&��M�n<�4�P�1Q��7R��)(Q�N�Iq,��� �|�v&�62���-�4���S�D-�׭�91m-&��P�"}��d02iL��j�"�/�/��1c�ϳ�>�f��x'�4�XL�]�fT"Bx���L��r�OH ��,8�)vSc^4�IX4v��"n�G�F�|�cM"�ڵN@e8P$�a:p Lk "y>y����Ijr�Ȩ�or-(9����z��a�6
�2B~�Ƃ�'�ڡS'�*�J�Fd�P�x0M�C�0��Ϡ�e
{�LeQ
�e!-8�a������y�m�}��zɈ5����z�ߨ�6LB�������D䬦�.�H�6�d�@�L��!3�RK�C�v&7��ȤS��u]���p(2iXK��b�'&�ߊN;Lh�y���%�1ۊ�������<a�ڻP,�U]$fl�J8L��ɤW j�,��S7�W@��&��`� ����z� -���w��MȉYU���}"
V&/F��1�ԅ��K�{�#�s}]���Ea�5�|�)Si% #3(��#�gb�٭of��H�3�{e���64+������B�"u"���N���\��yE���c:�,5�/
<D�
4�d�a��4u�[$N��׃��)���d��+�Bx0l�v�)�(oI[�*5˄�$*-)+%�2v7T����12���ji��y���*���N)ʰ�d����ٰ�w���W��}��D5X���Ȅ�w��]2�ScdbH�k���2��>�10^�`�L߫�P��^���{0��WM<��/�u�3b/�F�iS��%�Db�9��	�Fiݺu��JSS�� ������ �\�]/D�4�{�8�ыI+5�    IDATi|⃇aZ���m�����~ �XS@�8����Fz������W�~�n�=����{턬���h���λ�V��v���໑w�k�-w��>tT#XQG��wa��6���/�?�?>�/zJR_$('P1��Wŗg\'_�e@T�`��M�}j���NY�����3��-��d-��nh{����Yx�V�/��q��S0>�����s�<�j� ��9�M���Zy��V��/KJn��z��4d�n�Rx���h����L@֨Jją�Ǟ[�u�P��b�>oC&,K/�̟��
��(��5��D@MG:e�&SR�� [/�I}���m��,j�!HIk'i�E��j�O<��Eihr���� ? �@\�g�	�~5��c�����x�>�A	z-T�HM�P��5��`���>��&���ȗo䘆�և�.yrH^�}c޶݃ɍ�<9���oh#�84Z��aF��L��7�m&S7T�6��iS���P�˔ԑi��#�4���.:[W�G]�;p�>;�u�Z�����a��>�W)ê��߻?��Ә>u2����p�n����F���\��6�����8�3G��z�j�Yيξ=��8p?���F�� �4�:����ۑw4�yٹ�^o�J5��x,�ş���!cg��6��S��
�QUNM�����3��~��l\s�1(�tA�5�f=���Exi��4�	W�p&�L�y@�x��-���¸�:,�p.v۩#���Ew��܄��f�}��8t�I�X|���?�s.Y(iÏ�0�q����lkJ&�|�\��p�>�㲹_CNwE)���p�y��/�D6c��E�c|��� l\��F����a�5!��<��2��R��a7X�Ը�b����&&�˕�O$�H7�	5xքſ�j�1o̭��}���%464�1�,��L]�����ȩ�`��"F�x�t�!��~� ���]��L���c-gο�]"��D���ӹ�m�vU6:�I,��VQ(�Ij���	��_L�H,m�� ���v�*XZ�r5D9p`9)�Up�K�1%O>k�8\t�I����Pf<N��J<��J��^��q��S�vo�����y��1�������� (o���ÿVw�3 7���YSp�9�#����S�S8�������Rx��U`j��\��8W��\��VLn�	�J�1���[�4;��^���R���Ο{4�b;Q���)߽Ͻ���2?<�[h:a�ȓn�w.[���?-)���?�1=��jh��w=��7���Ͳ�{��ػ��W�AUK��gW����k�o�~'N��B/���S����s��}8`����S�F&,	պ���s/�O=�"fL��y���Y-y���T��/���������T
e�*��tv���H7�`�~�#̈�i����e��$��ȿG���=`��%������k��o�`r�/��o�H�Dj�U�Cz�,�����:���qli�ˤS���FDv��76HG�G�XɵWai��p�a�����)����w�1	�s2�,W
�H5�����X���E9��5��ۛ�7ᶻ�����&^�Q_����{��`�<��p��#�S8`��q��߂�d6|�5p����g_DC>�%��-��|A*�����n��uM(U|��@
ľLB�`ɤ�P�>ω�F,U��6?��D�^Dz�b���g]��W�a�\r�\L�+� ӄ�^�|�Y��Y|����n�P-�#�،[�{\}ݭҁ?�o�=�팠R����#ϼ �A����S�;�W�~O�Ƒ�8]%�����=VX��Y�u������s/aڔ���9gb֤&����.��j����`�Q�9Oځ�Hg�Pv9c���#!-ʱ���<�Z"��A�y)$_P^dL�"��iط�go�`r�o�7Ͻ��N���8��B<�)�J�!GE�0���q��N�o�>JzAL�땀#���TچE����tW�$�y���Y�&㸣�����R�f��z�����ј9��[B:_���� ~��{`�)|��������Ъdrux�ŕ�l��X�a�|��/ ���Χ0�w�|���u��{$v�6I���,�����s-��SYT-�55CE�aqV��h"�����V����8��#�G��}���b��z=fL�����jN	{�����<�L&�K�s:�&-�jï��+~����5|����߹'��>X�,z�\��薃��|�SEԻN�.;��_fΘ����u�:Udٸ|��X�ֆ�\
'w&4��)Н:,��f,�)��,�]_�.��������r0bj��nȑDg���zF�Yj�F� &���\y�׶ō�z�s,2y=����w���w���+�gC&2M02���ÑA$��Y�fItBT"�¦C�Nhdv�i'���m(�*Hg2"��׳�+����Iz~��x�;�Fc.��>�6�
��
��{:�L��@��J������t�\��r�Fc6�T���-Q��Ή��ǚ���6"4���hj��������wҒ2����JE8�<���B�G���y��(Td#�!��Z�e�d�)�Y��e$�Q"��eD���RR\��x��#3�^7�FfG�e�-!Ź�Q�r��zK>����>��Yw�!��PFhZ�hUd��ǩ9�[X�&9ͅ��ʺt��P�zr>z�^�MK��3�0%Y�-<��j,��'��,BFa1����$&`d�2Ek�歒YW�� ��Ȅ�M�b�H�TF+�lll�X�d��-9��Ln��Ɠ\�Ej��kD#�?�UF-��g�>��k�D���3�pc��O^/sG|?V���y�aR5֫(J(i�n?�������_R�XdKGT�E�`#)�i�L6��(E�Kg��J#��C�⡯�M��LRdoC� Ͳa��!��,4#0���Q�,dr9�u�2��}�~���G���B������@����c3Y�1�����I&�ɪ.��C�(�n��M��؍��=�iy�7�Ľ�K��ЊSF$F���F����I�ɒ�4h�BUO!480,�W�C����`�A_Ń�iP2���b�OтS&I
�8�$dD���Dd�	�υD�������;����@O� &JNG���q1=HG\Q5�WNd��L��<~��W�6�"�10�Ӻ�f��������M0��'ʈ�6"�B�v쮨�",���-��0��]Rh�6m��F֭k�v=O
�J�Qɯ��*�PE+N��G��=����y��b	��yT�:���%�dT9��u���Ϫ�I+M�j�l:��
Ӭ.�E��
��u�
�:�KY�|���ʙ�;7�s�*�x���o�0l�ԣPtL�ai,�)-!�Y����d�H3xp�J��q��Ҧ�d���j*}F@a��͟Q�J�
��>�6\ÁW%��Q�vP)�Ic%#	?2��^%����nbXi��*2"9`z��K@����a����r7���-��v�WUJ�q$����x�Mh-�����{e���B����-}h:+i���W��	F��Bg����h-���Ɏ[r�;�02!�4�� f�����|ʐfB��$�|^(�����N�2Uh��]��ǨEM5d�E�b�p�^|�S������BW�4LF��0
`#u�|}3*�q��0��i|��یT"�t,�# o_S*���	��T�J=�Q�h��8�A`q�6IW������2 �2aF�4N�������Ȏu��*�E�!mAh��#�2iRL1��32R��<O_�w��<	��}(<o�@#c��χ�h�C6�9�T!���*��YI�В�!�)܅R��A٭��La�Q����J�jd��:�
��q����0���k�����IpKE&�?Ĳ R���r^t&d$(W�0�R���0đ`4��$�<��gOXr������5&[bZw���P`���74"��C�XF��ϚI �R�k�Ǐ�t�	*ԹZ�z5��Cz@�#ί'��[-B�ڭ�d�i(w���[Urz̙|���b�aJT��N,Ee�趀	�mi'@����0Z ���sR�f
���:�!�,H�ǃ��J˄R��*�Ċ������^:sB�tՎǦ4��L8؋��an�W@+F<�Br��a�)RƗ����Q��Ms�s(��vTKչ��xR�IY�.yW��)4�M'�b�"둫ˣT�$��e9֔���1�E�)V"X��*8�ľ�CG��ނ�eU#+Q�3����$ť�9�� ���~F ��Qb"[��d��#.��dM��Rϭ�	J8p��%��`�x�������:k��dǃ��g�C��tu�k�l����%Tz�������m�^A���ѩ4�$����SB7�z��T~#���1�02Ѭ�꼯�"Coe���� i����E�����l��0VZRK��I0 �Y�" �T!î����n���Y���P�*�Yzn�vk��JR3doP(;#�)�k8s�W�h��";IW�"JBI� !g���j�}���/�'!�H� ��!�<C���D��^8����|�X�b=�M���ZSl岒�	���W�mq�+�#��	��b�LjX��Ɇ��E����,j5��`�L�WV�m�`:��dHg��1tI�q�Sw>L'��M>T������y&��iqLvt���w(0��τ��wu���dS��{���!��D�(�%r H�h�&&@�,fB�3�qjD�����O�����ʆ5�eh6_����1n�D��S��^?=\��	�u��ْj��+�-�S1q~^RGb�Y�tv}+�#jP�+�5�������K�k���4v��	�"Z2#����Tʭ��{2j���#��uS���?E:+���L��kT��!Q�`ĸ.���DD��"?3�z�DB�f���)SedйU�>�z���	�LD��u�P�q��[�R`��XK�0%hH� xs}d�L\H��qPdS@��48vZjl|-kaQ� 5)��v0YtͲﴷ��;��AJ�
l�`��G�Ͻ��U�W`��_z��Z���#�bŕɉ���P���I#�ʊ'��H�aY	���� �������O�����sLhwh$��g4�k�d���ϡOF�ƭ®R�1�87�1���*:�䊚��fL�����ԃ�	��؃�M14%���!t�8"���iw�[�L�5M�"�g��ڒ c�����8�0L��LY$74L)�<�y��F$�X�HK�ۀp&;�a8ӝTm�>��o�J��O�kƁe�Ft�:.\t�D&���H�祾c0��d?���Z	�
^��)Z.��]���@1�a�)�"��źYP�j���\yڨ�SY�hٹ��m��10������n�qR�}I�p��M��l6����qKd$e3�h�>�T*#i��h�;&��r�, p��_�a���O���9n�Z�Ua�@���fq�!��L�/���il�i�]��1H�p����;�R�U�ʨ��)�/�|5��u�m�-%|VZ9�@
�_"���ĺ���s�P�D���=uH*j�{�
\+6.��!8���z�����T
�R�a�"�(�= }�=X��%)~O�0'O����G��,@+?���hkm� ���u��(G������h��YB�����(c�W�m����/l1e
ܱa���Ee�j(�x�
�6��9ݒ�5��)>3�`��S9�����10�
Ln����}������9�w<��]�&oH�d�(�\�װ�$Z���];���'�ID"��1#̀�[0¢�	�^��۔�m�J�����` {'�ʊ�u��Q�� �Đ�.kvn�V��z�~���
��l;0h�֕�)�\�6!A��P�G���t��l�@���$�l	& @���+dE�����r�L�����wtI���.��lN�����	�|�����v1�xt9����M���g��/�u�����Q����y�Y�^R|� X�q��Y�p�⛰�߀��E._�dh�SP�o�Z��瞓�gTI�3� �"�|��2f�YS1m�d<��
�\�-&a��YR+y򩿣�,a��E0�o�NK��cs-Z����ֶ���`r{o��C�X[��*i����떡45ԣ�X��1i����^�f�����UjKy�*�n��&�L���{q�^3P�\�5���rL�:�pJR���`R��#�ĥ��Dy�C�d 2I��r1�:�$2�MR�/�˥�#�YT�'�vĬ�D"���-�ႊ;���=%�.ZgR�!V�^�
�Z�������4,Z�k[;���o��W�
�	�}]�[�X�@ՓO>�yg���p?�L� ��AGW7��Ʒqҷ���:��aF�z��gLlS�LL6T�K�݆��������B1&���7>>����K�{.��6�u���w�}��3�C�ᴳ�����໧�#޽/n�ɃX�x9� �~��(��o�:ݥP:�yխ���gOZrϨz\zV[[��c`2&;��r�m�e#/g_�l��_TY���]{Wi�Yx��UdӲV���'3�I�M�����O�vE!�Iu����q؞�P��E U�>��a��J�2+\��;S��՟�l���ʚ�pَW�畛���z�j���M�F��V�;���z;8�@<�������?>�����oiS�j�JOO>�я�w���H�<��Bl�җ�$���="�͙3������]���'���C��ۋY3������ N:�$d����8�ēp���D���g�F�ꪫ�Gŏ�t�R~�;����b�'��u��a�bR��m@{E��K~��"++��B�N*'`��p�W>�������_���>�]fO�w��,���0��$����>��9W�~7��O�{�d�p��@9�\��aZ$f�r�־3Z��s�(�3Y����ֶ��dLv809u�m�%3��5����N���Dj�	�
�J9��D#�� �MlDC���|�w?U�`�#S#ҋ��p�'|�0��,:�%V�xc�`r���p ������6(�|"��mI�殻�Bss3�}�YL�2E���?�q�{�8�3p�m��G��?�a5���W�u~�ay�̙3���{���`���x����}M���#~�U����W}���w܁q�������ʕ+q�1���y�,��3YGa���&|�|��/�Lr����'�Akk�oJ����j/�x鏱��!��*%Iv���xp�2>x���T�{��ۿ�ń�F��%d����圿��}��γ�zp����FG}������uw��z3|+�/#�W�����w/8c��/\zF[[����d�ݫo�o���\��$�	�������8���$�-LF�Lx` H��zt���W��
�^	�ˆ8�{�K!~���W��?(�.]꾏�zH�<�J��w�����G?���~���ǑG)���Ӆ��׿D��#���wމ}��mmm���'���G��o�{�7v�yg��� �P�f�]v���g>#ש��Gu^x�i.�^��.�T�ۺ�K~�c�v���X���U<��sX�~�F�dU��fi�31�%��
�2���9{NkƃY��^�a�#߿���5�����?�{�~�����SOcFS����\n��/�6��3��B�}�7/���y�nl�E�Noom�pLފ&}�ӎ&�o�-Yy�j��(v��"���|�Jh��c��ɄD5ʝT��)��Kd"@2�n�l��L�����y����C"F4�4����J��k���Q(�ƾT*ᓟ�����/���������ZX˗/����[n�p v�}wջ������'>!���o��~��8��n�Z"wBi7|�|��D�E7�32!�p�$��To=�4��G���}1:���Ӂ���
�3g�x����®�f��c>%�鬫n��Vqܧ?�C~��v7���_���-8��K�cɭ?����D&lִ#�Lo��ޫ���n���͋.h'0T    IDAT����~������^ߵC�ɷ�Rx҂�XG�Tq,M��]�_��T�ZD�2P��A]c|���)�g�G��R�.��T�"E�Gd�F&4�ITP�;7?=pbF4�..��1�D�rbڊ'�����u������D���u�Y�Y]]]���`�t�K/�$����]wŁ���O �C��R�u����'�(�1c����XX�f5���#q��"e��L�0���ͦ�^��Q5ӒJc**��"�ρdG~����òk����o�m|�����/�S������Di.��y9��y�y̑rlg]�#lЛ��ց�=g��꾫���h3.�����������h�r[�x�{0��G�O�얞�Q/u�/$����2(��bB��I�vBg���+W��.�J�_�������?^�I�"���G@���gol`2<�%ʺ��!��e�$9���%J!@���<��|=�����/)�a��� �G"A�ߓ�̼y��|�z���X����������&!D�=;�,X��\��ٶ������կ���!50m�4�{jS5�[��d�3Ԉ����VT{Z���쑔ObA\+/�kZR\��ڂ!�6�f�EG�h@gO/�J7&4� 9����
-;�a�8�=��̿w���ܺ����K-;����c`�Ư�h��L����u��+��T]:�K����0g�zl�V���i�:^�u7܈��߂��(|3���2�h(�*as��|b�֒zQM�$1�4�|N�NGI�� �Ț$ A0H����A�c�*Q��}�"�Bp`
���E��}	H%�l~A�����G��^Ȥs99S���̶�.���T��V��	���y3B�mC�k҆��u)��FJi���"�_M7�@h��	H��q��`�e��2�Y�¯��~2B+K���i㮼w��'�62&�튽9ǻC�	%څ���%�J�}��8������<Q(�_��ј2�g�=�^� 7�v'~r��7�H��0Q�^]�*KG���[�Oj%IZ+�$啀K ��(�h���E���hV�����Nc����$�3�7*I���x�:�(��@�%�+�Z�dx�#O<�	6׭X�!JՋ�&
]h��Pn}�_A�Ѡ��A)��R��MJ�����ʄ
{�;J�����Z$O�=z�6%[4�1���{�1��d�¥����_<��9Fz�|�v&�u�ŷt32�Wf�D(�[)p��_��3&�yg@7<s�)�u�� 7��[n�o��8��K��֌L��j��5�4�f�"�t�S�qX��.�&��ӳg4@��A�	ǟ��S��j6# ��?��7m�*����X���B����N"��p�����b}��2ʚ�{�l� +V��켬��赢Ҿ\�T[��!�҂�>��#�36�F���,�]9�+�Ibg}�3f�tT,���?�����4עE�Nnom����i�˨��
L�w�;B��)�~xхX��Cy�^��z*>�ѽp�i�����	8@O��C���<�cbD�5�C9D�:���iz��[�H�9��=i��=y~.�Ej�o�לs�98�Ӷ�MRY	&��/�1�q����D�1�F7ɺ�,ˊ_�AX|�ܽ��7��Ҭj��L�de=RA�vx�/�
]�~'Jq���l��]�2�.�X"eC��1=����y:�f�<���L���~2�mp��V݈c�UV`� ����]2��:ʥ��"��rljh���P*W��[R	ݢ�s�㝇๗V⅕k�ojA��0�FQҼ�R]�P�E�u4-��'����� Bf�-�ۗ^z)~��_�?��?������O>Y�誫�#��#�J��f!����Rp�xH �ڏ�V�P|�V��\x�C��kS^I$��Gug�J�Ɯ��dd�P�7ڴد:���r�~4x&lZ4#�Vcx������Ǒ�$Tf�C1�(0)���h����(�g�ͣL/\���K�"��}�����a��b�I�Aǿ���r����6���]�U�=;M$�dPQL`��5�n�״�3FL�,"("I�"�Uל��	�⊒�iR�J��[��Q\��)��������{��{�9���v)S��'Sѐ��`K]2�29qz-m��i�Vц<ȊV�`��u	&�).�X����SO	=��h�*��`��Hu����/ C ��O?���,�ye����|�A����ￏs�=��~z��du5U�PQ�J���\!;Lz��50�uҴL;X�&�� �����
�/5xM:�	�t�^=�r�$��B��|�,��#��´�4!���GH�(��ӣHڭ`���U�tm5���49j�0iZ������	�<���`�	#�A��x.����<��sw�>0a�7���w0u�T�5$�yS�IGC�W��:��ݮ,��\-t�42�	b�]���={�(���>��o[9>��^s�5��;�*K��f�m�}��G�����J�8mHX��۷/���ZZ�pa&���W�<X�QͭE�_�ruSr�c&��"ЦE�?���D}�A:D��Zۯ����NeV�8����I��+L�^}(t��ѧ���`�wW��֪q!�����"HZ-����� `�Ε�^qi���l �bΒ�{���������J�k0(.<��ET$;����u/��zKh�!V�C��E+���D�s.��J��Ih�.�\�i�B�-�����NY�~�a����SN9�v��ѠA�D�G���8�P�w�ᇋ��i#F'�]v����[nUy1�/��R�)���r����-Z���Dף(ļ&�}��$�pO>��|։�~��IfdF�ɳ�?C�����n]:K?x;��Y5&6r����z��g�ԫ0a�za2�p�0�G�(�6?��wE�`��t���L&<�t� &�+6�L�9��߹�=�<��{��F<��v*��Kt����)��5N
Az��Ҵ\��s�y�9�й^~'��l:̒J�]���9�q�_�F��0޸8�:ɼy�p�	'Ḧ́B�w�}WD~,���T����/�Z����q��АQ�M�P+���_~9�;�8Y��y�H�}�Y\p�"Fl׮�!Y��+��#��#GJ����J$B`��yG}� �E]$`��d������s��gS����p�����c�ɏ٩̮�+�h���q�^2%n���?��y22���\����Z@��$�^9^r4�02��|��O�aooz��ݣ�z��j&Ŝ-M�ܿ0�p�S˙撞{�;0mK�d�R$� [o�	�m�9�o�G|������>��~�*E:0���,t&-��QT�_��e� O�/�3�#�'�(#���Rh�H�^ڰ�
̝:_���u�0��Jhw�T��4mi=�Ɉe	��\��y0%u��W@�3���.��0�b��(��M	tL�8	(={��`
�#�<��C�������������{�Ao��)�`[��d<fד�G���ѕ���o9l_E&a���d��D�����tQ̧�\��o�q���Ȥ�n-
�>�ˆ�>����l �bΒ�{���&�#$7�j�z(��s�͹�k�X��͙�Zf,Z�H���;.��{:��	-����eds�I�������ݖ�▫����_��o����{_��ivY0���W���#QI����̐����Y��U���N����8�r}��71k�,Y�Y`'�����!1SV"�3 5�]v�E\Ħ}1U"�믿^ �e�J�����[��//.�0�Ej.�Y<Xc������h����g���� �ϧ|����[o����c�Z֐�ʻ�~0�V|9m:ƍ����Ey)\hkЙ���L����5��P���"p���sR��Ε��j<�����$��ZI��R;1� }�T�izs5�ȄcOͻ���1d������[H�!Y$|TĴ$g4Z�s�둪��e�W9�ڂI�N�8ۛ7�O�*�$�U�Ӱ�6�9`���H���s@�E�G�����/O�BN�m���!b��C�2lյ=Λ�Y�PR�
�-[���F�#	L��;|7{.*Z��v�28�`����k&l⤌�h(T���@�D>zV�v�ߩA!��O�D�L�DW-�K/���v�	��Hos>��9k0o���ߙf��.�䲢BҐ�>��#m�	�63��0k<��#)��(�w��PX|�a$�>L����������/
ib���ƶު��?�ct2y�W?����HBz�02I���T}�R�� -��Y3�>8��C�JFnH.�oCP��l�-J2�z��H���?١s��/�l�F��L
��nԞ�+�	b#9���L�(��;r>ou�.�d,���%�(&$/S�#��!kR��2�r�|�Ld�-6�\8���)�L|�r�$�JiG�cŒ���&pŅ�_�K�Ԡ��54;&i	��0x���o�el@CGi�[v|)�֦9�Js,*�0;��˚O�Ypg�w�Gs�,�,�s���������;�<T�w�%}���?��O��k�h�H'�k���C���$��8@�`���ثW/����?L?�8�iQO�a��Z#��v�I42�Ȭ�� ���W_C�N]�D�z����7��u&�0�V+*��b�V�	�wj1��QW�_`:�k�K-�J<���¦q
p�"�)�:Ԧ�4�F�V75�?
����#F&�I0���e�>��`�b{:���l�1KG�q�=�l�ec���Gx��7�hir��d>��d]��D&*Sв�`�B3,���B��b3�Wd?�q�vX�f����f���D�a|.��{޹Ro�"����H��_~}����4w��Qa�~��/Zl�5���a����'�RëiX�6�xr�b�jg(��(�阶J���|���!�F�$E�0\l߱���jz�L�+�p<��F*|�p��s�p�B�v1��ƅ������|�O�5��a�c�Mh_�Km��I!��u�K�."��E��a�) ��7j�<Gs�x�K\?`0-۠�bE;vig��|��f��,��"&Fi�=���q?~g���Y@��dȐ!:t(n���m��J������?�Q����=2��쩡��y/X������*z�D��(o05դ-�\�'6��0�`���Qd��P���D�X���%
���oжM{TV��@\��ad��v*�0��i�z��`�kv��b���<��-�L8�H�͜����X>�44�RdI����^����A�k��a�����r�ҹ?��jj�ك��3�}|M�,�M����9�&,-��Z��w�����T/Y��Ӿ��/�����De+d� �^yw���p���HR&��Ua4�c�,(���?�R��A5������ӧc���8��3��㏉�F��<�4��`񝩢}��K�T��b���K//��-�L8)��So�>?���M����5	?[�2��� ��&��3�:�/.��ra{Q�N�"��u�XCs��I�Ȥ���=w��`��!͍�ci�´A��;�O����Y���@�[U�)�;Ｓ��7ݴ�ʹUh�8/�,�4{0y�Տ6�pȓ�L�y+��/��k��.�1���t9�ل�%M��7�!�E1���А�`DbR�k&���0ᵶ�`�	�#Ts�`���0#�����?KZ��u��N���.<�h������b�(JKKe�w�������X�0` �?��
�B�\e��*��"	'$��ԣL�8QĉLpb�=Z"2���"�p�</��?�>�/�u��0��iE~i���hd�\����xT}{�E����`��NJ���o�6o{�W���M���n-�!� ��%��<=\i�-yRV�q�������IQ��[� ���k&�_�x��?��LLS���m�"�{Y�*�`�.�P���	��C`EA�rY����������a�=O�,x��q*ԉ��4W!�M6U?Q���Yd�k��D���-Q�[p�-Rl�bK�-�0�L�F6��;#3��z��&Tc��\p�EEܷ��nl�ްq-����5���9���N�?�Fԕx�Ō�Rgr��7�OA���$�g��0-|>���� �!2!�����Q��5|�^;�wL��<�c��4��2cU�ސ<X��ӫ!�-n�n�}��l���Zd}��=�<������x�;��E�u�A6��"<��1ͅ۰1?�i@�����N����e�gDK+��:��3�әW����ֶ �:aӥ�V��(>d���s��!X0u���S*;�(촞g���>-��SaTȨ�0���̸����;F����}P��8�R��ʫ>�*/��捛Z�nW���Tt7�}F�&U��!�H��4��O����f+\y�?q�!�a�]vZ	&?Og��4W �1�M�!Nh������OR��K�d�]cί�������TM�P��������MuZ� +�b`�s�I%��Ex�_-˔Z	�^xS�Nr#�ƽy������L�YS���j���X�I���^PEә����mʬ��"l[l�kV,���ݷ�A�_�^�6Ơ[o�H��F]���j�|�P���/�f�^K�;0�ZR��0r��`+�����9JH�o.��N�0U�0��`���f=7��A��'���}5��}�ay��0��I�X��,kڱ�=�녓�0�P��X��0}E*1�g��p"���������Ŭy�������bÚI�^_ٶ��,�7Ns5U6Ws5��f���'f�>Zm���S1��2}�L�s��f�۴i�t:+��SO=;�'	X����ו�oVl0a���d\�,w5љL�3ɹ��2��_��[����`B����mb�m����7^y1�<�X�����ۆ��"<l4�z���ƻ��%��2��cx�N�͵���cUC���i
p���J^���5�ȣ��]=�T�Ҳ��:u�$��&�{��Y��s����n���������I!�z��kT`�I�W@�辊�����hpb6�G�y�;$' �h<��y?TўZ���9��ZdR�i[����aG"k�g�fj�Fo.Iӄz�ƑɚD��Eg�\��1��c��,���	���Ɣ��E�'�ݶm{��)���gj��;F(=��l�hg�9���>a}_��,6��vs*����	[�p�(Zdr�Kv���h���Ej��ԑl�C�%1�J\s�%�ѥ���F�����c�}�<��^�-[�sWU��'��NE��U����7�|#4^��)�c��E�������n�C�%o����.�/
s���WT�����)�d���g��}�`.�*}U��*��P�^�5���q�RX�
e5~~c%������dB0��Tш%��02��~&���L�����I��(�Z.��9Gx��ζjr���p�p��y�(�㒩��&(�#�8B6v$�4�����_�7[_`�vTקL�͜'
x��XA�F,����}����Ú�.��z�Kp�I{!S��O>��;Μ���l�g^x��#�+���V���%Ē4�F�ª#�]��ֶ _H,d|���B�Z�9h�B��Y$��cS�x$Jbb�������o�}�첨��ˇ~ 7�|����e2�������Q͖[n)���Lk��Y���j�����^_|�ئ(;��ԸPu�ȃ���7�\Xj�鑪��v����A��\�7�����d�1��I�曯c��0[Rc=7�$_�mة4��lשŰ�F]�����}���U/^<���L�&N�ZM��ذa�$��[&L�f
�F�Ls��H0Q:1������|��dN�"���������b�X���9�&Ls1���dICFj&S���;����}哎���\�	���N*����%����H�X�����o�[o��͜x��7��>#Z�2�Y3���*(Q�L����c���\��S���J#.�,>s1��'�1�K�/���x���%�#����q���^%;(>�����C�    IDAT�);��Z��*�T<7������?�ԭ�ܤ��o��?\ԩ!��V.�t	f���d�+yn�h���%͙5~�@r�H��X��D[}2�H���X��
c��'�]v�Qjc�YD�k�3a^�{�S��4Wa>������~������G^q����k�~�L�L�8A� �_��<(L����M�)�q���a��`z��F�׿�%ta���۲�'��~G������ ��D�	k&z$òe��ZP����?�p���L�̴��ںR�(�ꨯ��ͻ�G�v��Hİ�.�������9D�Z@��u�'�;��d�=�ZP�����r�*�C�!wCT�S[�0�B�`��ǉ����	�o�&���9��L��{oY�I8p�������Κ�J��kP,vmdJ��Ov�Opcd�[|W`�IÉG�n�F�R�Uƃ��\!C�;@R�)��ޅ���9�,! �54�$rw��qrRr�з��B>��?J�S�jztÒ�ɔ/�� h@��5�R;υ��4���+�j�cM`��0��Q����x����F�����Q��.��s��*�)#xn�8F�=��/�b!А����q�Z�L֬3�F�	 l.���\ i.׌��� QZ&`�H��`B�&2~��k���%8��cq�c��XV��-ڣ�F1�0^y�]D��!�`������_i���T��Z�u�3���S���A��~XK!��3�:�6������|3��������?�R��駟*��]�|9ڵ���b����Z"����Y�	N*'�~*j��kfZ��<#2ʨ�g�����eҜip"r��X�$������A@�)1�Ԍ3Fޏ'�����#$]�[�h��>8=O6n΃a[�l�*���'tFI%��n�g��{��R�� �x�mo«E��t��8z$�EZ�x�h!���3��%x<GAWF6�Jڭa���(g�z��R1�W7�4Ws��2(9�f�˃�w
~9�8f���8W�F*��z>�ұ|gZ�`�9�y�������1�a���\�����<"p=ei��BV����d�������XQ['@�5�(`��s6�d����)�X����k�z͙��������#%p�c�=�@��GࢋoĔ�5�#!�6`�#���~��~݁�/�B��T8_X�Q�*�)ܜ,�-���|��JJJ���D!�p'Ǩ�=W5�L}�}Y��G����6F�.]�ɹ�>�,!\s�������LP�V�st�[���q�����`pn��fqR�ҵ�|ϕ�ea}��t1񋯱hт|?wO���D�3��1�·)�KҠ	Á���S[�#;��������_�C��������ayM���N8��������W�D����s��jF��j�Jd�RI�^;w����6��X�L
	��a�q�m�	x02aZYR�������9O�Yc
��=�A�d��l�T��8�Ɇ���
���F�D���4��ɐ�K.��,\�B6~�M����]���A��x�D�kQ�$�Sɭ�*Y�|)JbQ�r�Qب<"����cY*��C�v	��R�]�����-7��E>������H�|�D&?~�s�q9�Q(�T�e�ziR\��ȈVL�����$#��N:I�uQP�T��;�A����`Μ9RG���q��#F.�u|��{o���G��W_�g�|*�v���፷ߒ�����^x�|6�s�6x�����<#F�D4�c�n]��NO��ŋ���4��#��!�ɼ��H҈�b�k��s��q�_����Qw����OF�-6�-��uu�׳X\�} ��y{�y�e���t��}�9�)��p;�'M8FT"ۘ[��{����k��}s�>h�D�L��a����ƣlNG@Q��|��hT��Ő�t��K*�
7e<'=��8R�^Ԧ���_�uk���>,n�}��n�����F��6�0�wL�5zy\3�d��O�⥹TdB0Ѽ�^DS\�}�6�W������g�A&�"���&]q�M�q�u����������xbs��v�� �K��^5�;+��*���."��<�Ҏ��d�5>_��>�)�ɩȇ$.�VĖ{8tʀ�{ЂPo[�xy+�'`8酖�gmgsYє�ᱫ&�Q����L�(��]��V�
�!i6'Y���,�cglީ>��3|��"������0��>=Ɍ������͉30��h[Y����p����㞐N���8&;u����k�����W�����L
i���0Q�H�#7C<(Vdt�"�t���qN��愴}��us��1��>���O�D�_�o�)k&�F �2�8�n\����.�$ۈ	�T'�Z�U�4b���͹¨bC1�����%�i��rYd����_��7��g)��L-��[w�ϼ�{z~i;d.��t�r5K�=� '��٤p��5��@��q�����SzE�U �D���wj�@Jo��/�~
�B(vXaM]G����l$SI��1���(�y9�FX��@q}�n����I��$����:SZlH�)^��x02	�\�NA�+�LԹ�-P�ha��\�Q��e8p�]�Ö����^�G��c��8��}�Lg1��7�[ۡ;6����X��?��Z��#����<�ĳ����32Ƀ�.=Z�zj�5M΂��=��Y�):�c��x�u��&�),M8�Uj�c�<�<�5S��8�<d]R4�yAf"���GdD�ȤPP��_�s�K0�Z�h��Ӏa�"4g]J�M,�K��3��>��5�������n���&�g�Д_eE��L/���D�c����t�j���r�DF��Kd'�Q���R;�G"W�7d
+��\��h�	����dR�.�x�QJ|>����E;��ru�� # 	�}��	�.4���G��;��`����r��q2�[q4�!��_dn���q��:K��ISW��j���I��b��c���2н,�t�vv�f<<�1���4tٸ-\�T/]�+�?�e+����?c��w���?��^z�6�~��E����<uF����$2ٱ{˻�=��g{����7W0il���M�95!�!0 X�cz�k	�%�	���#|-�u;\�w6�� %^9;�=9�Թ��w�>Ϸ.����d���9�T�`��t�`�ZG}]U�됄�o/�Ҝ-����h
x�L��L,��䮂 ���m+��2�/&OBΈ��&�J�?p2ؾצ�Z�f��oI*FF�����5�������@�q%��8b�H6U��℠��ܡ�9�&wh��0�̚�]x�ǹ#���'���i~��3ψ�=��B=���OF���@�z��#�N�����iS�q�8���Q����;�Ʉ���ဃ�k����CK�;�t&�O?�����'ow�#�q���|�fb�l�<�̭��X������f�nA6�c��+�=r/�>�!<���r�M1�ʾX�_���#�w���)GⰃ��/}�{|�t�뮾K�,ǍoC5�MF��E�k� &�A����n<IE���NZ>����0���p��0�E�<I$� 鄯g1�s��N�\���L��"`HԦ��ck�ܲ��3&���/�-DPZ&`�xq5L�^`�
dl��������#n��t߬'��G���"bj9�:������+� Z�N
�!ܙ�"�3��ݥ�gӺ�LT��Q'U,�sWEaA��x	��b���c��3��O���Y�N���![��C]Y��ؤ�4a���C#S�9�+��Bޗ6��T|���Fy���.���v������ݷb���˭��O�R��N�^�����cO8�&M£�m�m��F+Ĩ�_4Ns�y6W�暵"���~H�Z4߁�ˢ�Fm`�E*�Ê��\�[u(�����E`�h���E�4�zy-��t�1j�aE2���!�WF&Q7������W�Y�ﺘ�l��y�
�)��4��
�]dx�zʃ��B@��8�E�}��+뇌:$�S�p��������b~o�>�ڂ	�Ԁ���Y�a�(G��&l;�L�E��z,�I����%JX1d2̚�ŵS�dHh��
�x.�ܹ����p��[��8��y8�ҫ�y9<v�xh�x����+ڇ������"^ӡ+6�oLx�*�D0 �]1�Xdd�?��r°�H�"����PaN����t@�(�bDF�O�w�L�c� yp"1�L�_�����hL�0}֩S��u��{?���k��ㄡ���;˹�1�0�L&��ͷ܄�5+0n�c����%2�rvT���)_������$��u�h9�9�,�l*��m��0��B�k&��.�N�\s�^�j2+cKhτI��H�����@`���to5���W�Q�I����\��0B�<a�CymQE Q�8'��U*W���3M�.��ƻꪫV����]�8c�'(1\�g��=+�n��.�w�s��/�`�DM2��Kj���E��	��A�V]3�&���A�G<9[��T�4��3�~о8���0����ݫ��x�H�����<<0�_��'���+C�I>2����(N��<�r��fR�8i�H�A\�w��R;)Z>�_.�6�oF)�j!���?�t>������[�LFLP+BJ����v�T�3O̮tLm1��a?# �������zy�Em&�6��bI�RT/X����&}��%�aۭ�Nu��g�C{���v�O&}��N;�z������T$Ea��/�3Q
xO\FC�I&sj}8v�P�e`�,��p�
���B��BvZ�H�D���"9��qr��Ib+	yM�;tos��.?}]/��>_s�5�7����b�N1-�/�(�`)0`��l/����%��)bF6��Xcd"*DC:-2��9�:-�g�G&1�u��GcB������x��#k&iWòL�O��Vx�kZROe�h5�B0ak+�S��f3�f��p��H���"��������L�[����)��T�+��Ԉ�$\�����T�(��H�mt(�(|L��������i.���LkQ=��{H:�gϞ�,g?�J�E��>�:(R�:����u�@IP�N��d��6�`��%��ǋ ���R�MϽ�<�M��^y%|ǃ���_?Ѣt��U@� �4�\ǌ��W�ǅ������ɔDAb�I�,R�u=_3Y,�CA���d�D&�ژ�I �d~��
��S�=�Fʰ	��-0�W�iN	y@�8q9:tS(�ϚI�1��촦�Ȍ�k�EUUU�5G��5}��2"�]�F�ĕ+��zn<�;w�QGɆ��p��`�3ӣe�W-�7�>F��$b�ͺB�/�(GM]��K�t-�e�\+�&Sf�A�}�"Q�F�Z�_6��Y�L�\�2+L&�jpDs�SRp�͈�V3Nط�$��d)�%�X)�fa���"x&b�v���L
�duCJ�a9�).$�(%:uZH0�'�`�!�"�(RYH��h���4U���+����(^d��I&�6�Lj��3��/���?>���t�2I_�6���/�}-�D��V�+��5|�HdG}4�67�t���g�yv�}9SW��0�<5�L�&-Q�60h�8̫��q��$0/x ��.����f��ȧN��Hҟ�jl2���l/����0�b6��˳"���ˈc�ԩ��ë́�3�W�Tb�`݄��	���G�ٗ�F0)�/��`T/0iSj#U��ax�^���E�$&�EYiB"�l���ڔ�����Po��K��`��I�`O'�=��R�߸u9zo�	Q��ƞ���&X jk�`Y��H�>"Z���(.l�B?�35Eο6F��Y�R�W��)J��lU�W�`��X���/:�da1uD���r���3�g^����gdA�zשHW�����4�|o2�x..�L��|<�ԒD`�sϽ���l�u�i�b�-zJa���g�>�?N8N�p��Gp��� �S�1C��ο ���!}L��'=�Nņ^R�C0�S�Ww_;m��h[e �J�E�y0	#��nGh�ALz��❗���g�o䉿��D9F(���1�q�,�	 ���o�k+�e�L
�\B���?�j!���)Z%LXZ����RR�aF����Ԥ�:)���,���L�3���,-����]�4WadB�"�q�d�LZ�7�?qnbs��[�h�=zT�Pq�C����`�+`r��/"_�#1��E��-�l�] �֠��c����a)��7g��Ce��ﾫ0�d�Щq����ߕ���R[����<`�yq5^D�Щ�S�_�&/T�����Rʧ���qaj��YZ� �9k6�v난�k��Q��z�����r�eD9��1qa�1Qχ���	`ږ�ɪ���}Y0Ji�F&sk}�Lh(��� /z�a���NG�����0�ӣݘ�Ｔɥ��{l���U�oi���+9�yF���G�D4ɚ�藂��x��Iy��2�,|�Vb%�FG����9~�� �`��r�x�12a��4X1c��s3<-zK�@��'v�m/�j��8�� j��p�x�ɥ���at�=��'�+0YX��$� p~���p�p��3�(,�'�@��Qקvi��ޗ���
A���tD�Mu�juY�}xd�:��+O�5��I�aE����{�敋����2YĢ1���O L�bM`�v�ʅ�S@v��N^O��4X!c���/��UV;��?���/��&�i.:���a��w^���\�S0)$�4�ƛ95o�4o���L�ܪ��9�s�X�T������:t�6ö��:)M���L�f�q����%21��+�3QSR�H|<Hc�����`Z�ԋx�7��_�XydK;!�(� +<h��P��|Vl��TTs���A�"�_��� T�U�U�����F�
m���V�+�V�Ha�^U�)T�a�`Za�v��CQ\8���iI� ��fX!��g�b��͊th� ¼��t&-�F-�O�}e�$�g��4�V &�L´�O����������eU-����`һ�Fw�r��MN?��1WUU��E&26m��Sm�����ߦ��5�IAͤ0�,Y�Y�&"���S��I�E ʚ��U����pr7�r�g��c������I�;���J��C�II�,]C��-1��Ѿ�ț���'H�ۨL/��_�Č�-��*0��J�3�������葋h�s(m�H�p��#+	�.�i�cbZ�z�?xR{Y'a-BM�g!�^�Rz��a�|�F��B0*��j�8S;�B~a]h�����˽H��q��
=��� �|�13XQ�6#�~���{�
�jX�K�sj�g��ϤZ4"���5љ,I<f����8=�%--t>3_	��Ta���*z��lZ�B*t]y��tX��Ȋ��`�Mڍ|�΋�����L~P�Λ�M��LP�X��z� ,��ܯ&#�琩�Eİ%I�2�l�l
��ی ��J��\���X�D�[��E&���a���?+m�#��TN:��"ͬ�V���B����ѪE�Y������f�BX%���u\���),�����W[3�!?��v�-��;K]��r+�n�fN��H=���7���̓�p��~�[�*@b�������_4�~�j�� ���_��Z�xM��}��-ȩ�V�EԶPa<l�8p�}p�q�c�������p��'�����? bƞ�l�?�`�r,��#��U����v�쬃tćӺ�G�r������H�0i�W!�K���=Q��i��<�9u9�f	X$��
.�$����X�����V ~b�-�!0WR�Cʸ-Q�����l'�m��{y�M�9�=w��d��[����:�O�_#�ȢI�N+�XV�yӧ@��"a��$Sa�2ܢ!VC&���DX��&��Y�ẍ́OWq�%�"�Ƀ�|ܵ��q3�f9���j�,�i-�\�t�#:t'	����X���̈4IJ;��[�.��8�    IDAT��a���٥�/`B���C�X)v�q�Q��}a&o��O?�X�}\��S�ի��(A���[!Ł��"c��{��]�x�O<��i�+dJ��KK��&Y���ː}��J~�!��"8�����FM�S�B���æ�����?~9zH}��6A������{��Ӑ�ӨK�Xڮ�f�R�N|�B�0I:-V�5$�X�
,Ά���u.<�&"���Z(@ ���� w	aG4��Vh�O��2���`�ٌ s�4V��v.��]W_T�{^�s�=��K��� &Ÿ�M��k�ե��|Is}�R�C,�#ېY�>�\D�!�H�S�D[-��
��E&���?3m�B�â*�T9��U�ͤ���Fe����eGQ��@��
b�'�^&ԥ�S���_��@�Dd/,(�Y1��.��@21�-O�������~�b?a9y�Jum������ϊ@�*sz�� HPD�
T�Sߡ�T<'�ԋ�ꁽ߷�f���-֐fM��E��P���l)��G�G�ZU��_�;C���.�ig��u58�Ŀ�ˤ���;`�W�x�'��sOF׭��+G���)�l5��E�}��v�^</p`i�M��U�	���5fI9�2ds��4�o��ԙ0�1#�60�@"R����,�x�51�@�9̐4yѢFӺ\�7����]��D���K�r����^���Xw�i��I�� /l��Qii�X��
u9������u2+��_L.�㱙i�Lz��=3"(�بeBwS�45558���Ѿcg\w�M��T �ٹ+5��5��X^g�#i.�)(C0�s��e������Cn��/�H���6
Y'Q5���48$�0ʢ�/A�V&�Y�X�F(6��"��>
��\�� B .�6Y�#�lT��	z=���'}�cN9�:v�.[l�{�����Ǟxf̟��/:Z*��>�J[`D�~8�信�V[�c�F.��42����2�}n_������LY�bk=}�X��J�����2,���`Rg�;4SY��"=7mQ�8t����i�>"�g�u�L���QѵP�����3X�g,k�.l�%׾8����ǽ_��1��1�UUU߲!2Y�w��k�`�Osy��&ԙ,^�o&}�2���*�0��� ��e�]ʯ&S����̬Q���ƴ���dRK�ґ�8�Z8�N<�t��}/�m6���.>a�}�Q�Ju��ȤĈ`ϽwME6���y����`�\�������QDH@am�jZ���q�ǔ�;#��;�8iʃ�~>�����zKx�@���	'���]�J����(�����3ΐv���4��G���z-۷��o���_|Çŧ���p,&Ϙ�eK�p��{�OC��7��3O���*�7/�HM*`!K���ܾ(�?�	�Cϴ铦�j�R8ºbmݗ�da�����1�NC`&�k)�<�a�~�!�.C]�WXgQ:�s��
#v*�W&i��) ��XV)4���=�]�������o �u}G����&�4K�U�(A:o��l�,�;j��Sʬ{��1����D"��i���}�/�2�㛍�R�R��IO\s�MR3�k%B	�`��+�>���ɚ���	�j$t[�\�M�z�9O<�$��O)����aEF�R�!Ҳ�O�J��J��>X:�� �y�Rئ'�Z����/������nb�v�r2��5���U��Bb#�޽{�۽��{�~�]�Z�m��v��=�P{����<��.����O�'�G��!	����S��I���2b�x�,L���o��7� �J��i��Dբ��9��`��L,�Lf����8"��x4)譒��]�3l
�����)lT��K[T*�\��FP2$���>R�	Go�3��&�.y����u��u�`R�;۴��s��
��c���!��S+����I�|�
�������]��J��	��#�h4�� ��,����L�����@g�>2q����ㄖ*���Ms��VjFW���M�8�|���?x��Xd' ��E��|Pb���I��ф��A�R�'0��m�ݤ�M�iӦ�62
a���ϖ���`RHI.�V&�J����)�f�����k�a���bi���\#���=����wƃ>	K�Ю�u�Z�����a¹��$�A}��8@�������\K`x��su݇&`b�F��j=x$_58�Aml/�s`g4ٸ-�Jt�,�A�dv���]}Ĵ�m'.�{3p�a	��1��E9�y�����}�-�?:d�-ż��8�0)�]m����`"��N�L�3q����@E��=p�Ix�'m0����L��DT,3���Ja���n���QC2-��x�(?��>� ���f���𼁼�����~�!��mfo��&1K�������ѣ��AC9F*�;w�ş�0{%�ɔ-A����"I�e��C9�25�z	�g4h�M6u'dR����v�P5���WᱶD�-����:Pt%�W&���c���ȋd��:7����F�:v�XH�}8���_N��EKa9��2����U���a,���N`�ʹ�%2χ��z��	�Ɂ�eC0Iסc����{J�m�F��\R3��L�H6R���T�w>�&6�t����5���q���{l �uy7�Ϲ�&�CДWc0Q5�Y�����b�z*�1�5����}/M���·f1�E�-T�*�|Wj
�n�-�>�8<���x��`X1�vT�OZ0�^Y�_Y��&�:jq�1�	�\��)��.��$�\KVDl��ڶPh�H���!�E�ԡ�[dc�ź��<�E
��
k)����#��KwS�Ja��SC{u"�u:B�]q=�}��2�����4�	���ƒ�E$}��1�ۮ@�.����/u �����`��*�X%rl~� ޲�$}��A,Ni��(�t,�:�s⦎t�r�W����(�uXu�����C��K�'�i��P/�8��\�� F'uZ4D�`���e�>8jT�csm �u:����&��##��?�������F"�'f���,��}.�eH�,�i�����O���w݃����!���P^ٚ%T)���%��h�ф�l�=�j0�%���hF�{gZ�Ju��Z�j%�ʹSV3g�S^��*�1�,W���	�6�)��g��
S]�d�������?��|:J
ty ���}w��ba���A�����m(�A��v�4��#���o0s�<��Ś��*[`����:v��i���>u�E��p���M�W��2,��x���0q�(�&`7,���b\{���i���ksa�������b	݋�V����5w>�r���F�}IS[M6�IS�����6{0as�K�=>;i�����#QI����uKѶ,���;�@L�z&j�YX��s?,Y7��6*m[YCQEw�c�����o�
x�Z�%`�۞����w<� n�9"SUl����_�W�32����Y4V��T�*RȂ;��$�_X|g�v��_(l��COE*��k����#�K�5y�����&Z&ü`�$d�0�J #��&�a�K#�f�� ӧ��w��I��kgO�Xi9$���{�j5i���9�͉{i��\��F�3���*�
�s�x���Q^�vj9�4���vf �����am�d�=��#������(������.�������{y������o�q�0�x���f�xqq�M��Ad�Yhn��B��%8t�=p���	Ӿ��e5ub����Ob�����^'�Y�	�\,��5�m���PN�h���B�EFQ�]�Jwe��:[��!�����e�K��9xm�����J���ƪ���aHX"ӈ�\1� �>^k"B�%����hB����%�s��4q*��.�k����疖a~��mc���zKt&�F7iF]5�>���5�-���V��$�6i>��6�:�h��7��3��%�l�u�1��[�)v
5NNdc,�{��-����l���tm���~�0Y�w�i��� L&v�7�!qm|��f����q�?���uu������S�[1d�6��'VT� ʛku_m�,�o.*z����;�K�N�E�i.��z�,���H�B2�F<NML�U��I�O%k,.��X,�zaHўY�5+�c�u�D�J~]D��Jq������Y��hy�9!����r]� �N	�LSx��f�Z:z� @"R���"��	y�T�.^��3�HM-�`�k>"%eX���(�g"�j4zuSHd��̿�]:��U0� 5ZK�zq&ޟAjrkXAZz3p��`�.P�ϑt�Sr4�tE~�f�VX�^��G`��b��M�f�L��⾾��كɘ&v�b�ó3y�"���v���>{쌾���Gއ�_{f4!������f4���zDc	|M�(T��\��F�,�(<�Ҋ�������F�.�b:#�� AQ!c��Q�Q�З��'>��V�I�8	|���Y�����W�,[�~<T�������+i{���h������Y<?�i���S`��Pe.�Z*�pQ����9���8��L��Mآ��I��MX$MД.�L��u�_ף��(�l݇UZ�Ů����Z�U
�0�����V�S��{u	P�%��k��c�3���,�x;�
��`��`��sP�/ qu.}�e����L=@��
�-q�-�ݨ�-O������k�~��=��ŋ�nڐ�Z�;ټ^�� ��#��&�+biH'S�����"b�h]Y
�k��]�xԆmG�(�D`�X^׀��� ��q���j��&�lVj&T��6�\)�Ld����^�.��-�-��L&���7�R��Ć|��9�us:�@@!����O�Ƙ&#�p������{����l�I�nr\���Yc0Q � K���{) R UpN ���*�l�K;�Nʶ���!G-��!j�H7$�%�K3�2�^XۇaR3��bJ�E���b�G��#XX��"��1h�:��58��>ؿ��Ro!|/�t�#n{j>��Í���/CI��� �ڡe�"�P��J,χ)�2Z,�{�ܛE��v������e�׭�G�{eu��7��:����T�Lx�N?��E�ɢ4O|���d��f]�#��W�G�4D���L\�� ���C1c�,��Që#4�s��`$\��b���3��{l���0��Z>��&�9���(��ˆe#�N���|eS&F#�IaD��e`�V�{��e��E��i�o�HV_/� �J	>��0Ѵ��̅�m�V���uK
�|��d��>_�Q���Q��i7Y�=�{�
k'
LD����h�w
��ߙ�o� '���*�3�����\I$"�e�2h�#�N�������d$ZəÄ�R�J�,]C]��E�La���H�][��.Kih��0�Jvr!�8l{�(wK�h�۟_�	�=Ԣ	+�V������{�z$�E�PQct�܆���^�=Y�q��!���>����c��^\u�0i�?�Z����.��C�l0EO�����u4T��Ђ����`�E;bZ�dS�N:���zo�	��	Z�l�A�o�ŗ�Ǣ%�qϽ��G����Be�6�9���*	?t��Λ��\���}���=�,A��:���!D`�rb&���%j�J+��f�lIU�~��&Hd�)�"lS�w+�v�T��X�Li���q�0�H�\N܄��� S�E!!�䵬� )�������n�r�I�2��F��$Z��� f�I����t���ܶ,_��%�s5�S���t��a��䄶M"D,�@�ÿ�6A4U۲�r��������}�=���vL�Xٺ���$�� ���V
��E�u��΍D\�=IF� k��Z/�#��YD����Zj)��I�|�v8���r�\�2�n}�;L��"k-���oq��;b�5H`�اp<02!�P�����C�h���{�n�g�Sw�hz`2j���U�l �u�7�S�0	购K놰g����
�L�τ=����0����s�E���4*+�d�Kׯ���'q�8�dTV��f[l�IS�bYm�}�!<�ؿ��ko@�lX��P�W�0	[��\�Y��n�pR8�ð�6=M/A�k�E�4�N�	v��4j#�8 A�0���Spw�#��� ���&���q
:����G�8��s�f�����D��Mĺ�痣��|l�;� �x��ĥ]{�G"�R�k?;����*x9W ��I ��{�(���e������0v���@.������y��:{����5!�%�K��M�׀ZRק���('K ��\|nDunEQ�Yr�a*�T�@C�C���m����:��"���>�yu9����eԃݰ��v�`�"��	��Ƹ��/��W������ԡS�[8gO��e!������s��I$�.�Fk,2�Ź7�Cd�>�:�ɉ�5����UWo �f� ��#L�x��!=3��g�����W>�x���sSf|'���8jWԠ$C6Y�Ҩ�q�Ͼ��{��ӎ�����^�ϹKV�"��n�J��*���>h�����Ұ�,���A�s�-s�W��-�+
긘Ӓ��`�J� ͻ�hV����<�E��
}lriD�]�`�*`FX�q�Kף����#+��>P� H�� y�j�h�mC�ؙ"�@�؂=�o�>��/��#<��:�	�)�\�����oQ`.�Ú��2J���,���sF`5����D}6?R͎JJ��fb��L*-�� .Sf�T�^��[d*L��KJ�|��.ŁL#������'ֲ�Y�H4#�D)��|�U�B6U]������5q�бp�r8$4xix��
�_p"�޴��R8��c����O��Y�v��j���s���=�#���Q̨��ٵ�xҜ����Xdn�ndd�{п�mz��Qco����b��Õ���w&��e���B�L�#�E��6��k�C&������{�³/�����I��MX'�!��I/N6)��\�]6n�m����[�����m�h�������OBZh���[tE��-��d��X�_~3[j1[o�	���
A.	�$�����C3c�Hk�]�G�_+�\�^z{jj�hY��}6G��\����YUr��|�Ў��$����#�lG���1?5A�c�8�۱'t'�@�P�x��˺(�t�}/����lH�����v��iQ�=��r�*vF�_�_�	�	M7�ˎۣc�R��,;��U�1a�T8���]:c��݁t��TM6�[�,���z�^;"nx��s5�<�����N��,֙J[��w&��Gt�6�Ѣx���`�7�إ0⺏ [��|�yأg-V$bX�n|�<����ʃ������;|�8f�� �+K���hQ̳I�-�[��ơ�]���5lX�����3j���U�o �����z`r��Υ�#�@d�p�d���OI�FÒ��(��K�n�l��\����L�EY����o�Ƃ�a����x݈��pY<�L����Z�(��l֡n��"��Y�,����7�{S���c���Ыc�nF���4#x�i���Ƒ�n���E����ܥ����H9v�nk�����	�-tJp���0wazv�7�:VD�kL|�]Qp/͚Xސ[ieO�WIԖ�|�ן��td��ǎ�j����p�y' ��a�J��w�h|��<���C��]K}�&ܒ�q�����[�"jx����s�rI��r<���u���{��߹�o��a�<�ƧS����k�Ӂ{��ӎ��Y!��o�fqv��PU�E�]1����2S��.�����8;�*�S{��uw:���P@��q>G��uPdQe@T @�m��}ܐEd�{K�o�����U�L�ǯ��[�U��ꞻ�{���C��q���e]Y_�,�S+���[���9k�
0	n����<|�{y���NH���
�    IDAT��u�}hǚ�,�ts&�Ň�~4�9�B�k%�ȾJ�3�b��
i	��\k��ԏ~վ#.��k�;���������������ςɞ_�}y�3`¦E��NLI�]����*���0����2җF����Ll,��C�4ݖ�E�񾤮\��I�u�c�\W}���[C�S�é�]�[�܀�Z�x��z`yp�5\��_�뾂vj┷��w�,��-��
n�o��ѫ������?O{�� `�XTp���ƽ��O��>��0׍��G�܅��[���?�%��b7|I-ٮ�ޞ9���(�S��|g���h�j��_�O��(b�B�����]�6��e�pљ��'oR��}�:�r�=��+�>�=t)Z�c�U|����g��1��v
�=�@U,����p�y	(��?���d�S�e6��M�l��3]��O�������|�:���&,�ۃ�9��RŇQ���.�?�߻��l����51Q�c9VM�w� _�5Dz���,��k2�WK&1�[�����p̲M(ilZT,�H�TX|gT"���^�O���,*}�_�� ]@���W����U+W_488p�,��kgnf��o
L�#fW2��!"�Co��ɱQ1*�d�h����Ԓ4�I�!�[T���KW	��x��R���r���
��cg�O*i�B/κ�r�����Tʸ���ᅇ-��������%���w�k6���W���\4�l�Y�Ư������c�����7��2Ы]��i���>�z��W.�(Vt$�	T��યވ+���=K0�����*��`�m��t��@��N��!݀u .z�[P�Z��H\ěμ����A�����?�>��a��^�Y܀o��7�7����w<eI/Z�0�u\��[p�g�,U����xɳ����v��u�e���s>��7��
��;e���}JRu���p٩�E���x��t�'p���+%\��,vC$~Z�_�_���p�
�L������n�x�8���v�����,$"̅�КDt�q�)�⹋7�����#�b$�-Q	�J
�����0�?�}�s��?��/_v�;g���[���k?104x�,����ݗ��W&����ϯ�̒��m�S�v�\�J3���H��!��P�^�@H�e�C�d{`B����k+�ˁ) b��11��?y�>���) I�Y�p��p���Hs�Eg��/�A4�s�����3\�����hx��o��;�ÛP��ŝ�o��οTRq�?�P|�Է�O��Ѻp���_����V]�!0���5�b��k��C\����ۻ?&Z!\Jń���M��c��ȚD���`�1 '���{��W�#�ԗY����.�F��Vx��N�<�3E#�����'���A��r�K���S�n�}����~$��7�/x���H��E���u���_��s�:'��p�Q�� �I�l5�C�.[�ӏ���C:5����X?<���.��u��7��Ub��_�]�G�Jm�h3t�'}9a�q�L�r�r��б]Ki�1Je�98u3��؈���%xޒAT���)�T��-GvYd�fH~��$����Q�wȊ��X��}̀���O��,��kgnf��o
L��)��"��IJ�����(�q�7e��MzLW�L(1��j*#�QZy{<lZ��%]%[XJ�M#���S2Q/p�h�G�0��P(��)�wW�t����m5��Jc�tu�b��Z���~�Z�5#¼�2��%L4[����S�ʐfB�D2�^5?�,.��!��N|�M�IV��͔T�(K�ǘ��Y|�塮�Ȑ�ZK�Z�$���T�����/����$������E�]���X/G8	w$���Iu0�9	a��#d��.Z��s/���::`�|�h���y�d��u�s�Dr����	tJ�^{����&P�T�"15r��RZ]dxyFƴ%8���ӷ�S_[yũ3{����_���O�wL�����[���k~tےs>�ٵ�L���&F'�IP��1j������]�
D��HՕ��,1'�('Q1���I��I8+E7��FQ�2d��A#��Ș.�wD�І�$^}5[��G`*r��H�5�����tdD-���ӊ�h���t�ic�ᧁVG��Sh��?�|����ٛ��Jh�i\���=��d��<!� ��x'���d�(��+qK~�P��eΆJi�T��.����eR	2� ����$9�~r=(0a.��T ac&��`L��"�s�����ڈB2)}5��)��R�Ґ�ʐ}NZ	��?�͟pȡ�]��K>��is]y�%C���}����}����ݶ��[��X4��`"FG��R�U����M�H�j��c�~E��#� ���,V��T���.�4T��Y����4�t�&����S��*A�l�Q,2!��,E�T��`?*es��P(�e#�s�RE��>L�����h`9(L�C&@B Fў��>+��?������~a��~s�`�9pB}��
��TE��32P��A8�ȉ#@;��P�A@IdԶe`X&�z�ֽ����"���yu=����iZ{-�<S��T#�-A���jd�dk(�k�H�9N�Xfz�ZY�F�~���'��О��gv��V^{����g�df�y_��_=�pl��}�!�f(�������j��P�I��y�~��u0QƉ�nn��z�=gIy1ߞQ��A�h��6�-So�3�9�5	 �&�t�,WdB��3*9`�B���v�B����%�&&�t����[#}��x��_��I���J������!#��`��ϣ�ܳ�q_ʫИ�����q��FL�i&B�i/NAԹJ����ѲR��
�XlI�d���ǇgxJ�_�T�j�j���V���`���T�S��Zt6iRݘJ��&�Ơ�,���$'jp��>��˹K#C�bٿ��[.���5���՗�2&�ڙ������n�s�i�|v��F�`BOXu�?<*��v�~ع���fF�;]?��?��)iǞ��R��73I5X4C����{��܇��R2�b�$@�a�h�j�27n�	�˖(=!��X)���D�q��Ѵ�LG�\Xd�����f�?�o���u
����>�d�I���&_�!��{�b�� �5I5�dg��Ɩ@I�^�I"@���l;�R"�,e�	4�kUi)#�ɨ���)�ר4����ԓc��LGM��ͣY�L��tlI?Z���gjQ�Y�j3����iBJ���J��e�ݟ�a�Uο���ϙ�[|�o���׮|�,����ݗ��W&W�x��3/��O�\�Л�;��t�G�AO�;�׿L@�f�T�T)�����Y�N�+-��)�,����I-��?���u��tap� ���(�{-������-̴5P���M���^�E���"F���R�5�.�T�����t��0r`�
&����ԏ&�r��^"�����y�"����`V�g���\Z!������2�L#q�:���~v���`���X���<�F��0a�x'%� fe5�lD�8*��c�4Q"���=8�W�92��R�	��y�t&x�DJ�_�DGl$�Z+Va��8ji���A0Y�����9&�������W&�o�ò��sv�	-Q,�O�靪>��Nd���S^SPB�jf��J��In�h�����%�4��ݔ��B�F��͒(SǋzbT�o�E�BU ްnzjUD?�008"C����-I�����Xk2b�y�)"�-��"&�����$��M�Z�듏+V�%�ŕ�%�k
i�%}E��s;����<�V�^F�SN���6#8���f"rFB�L9�^���3�|�cЙ���� �x��wn%�ǧΝ�S8*��f����ɇ}q��4�j*v��OBE&F�@��k�ZGS8l��Y0y��"
'Zlknϛ��->+�7&Eآ��b�2��������	$�u��%0ɢɝw$��H�Y�]�+B�W�.�'��,�k��"׶�P=��`�<ʰl^�ղ��ZUb����ò��9V-�0�y���
�MC�����*+/��#3�$�(�gU;����ԗS@Ƥ�/�<���"�Z�5%+MƕP�9?��4R���D�N0��;�hx)�����ddl��f�0�����s��`�"r0Q�Ǻ�*��,1QA`�Fj�A��F�"�~�!$a(�6*�Ƽ������+�0AE�pȢ��?Xy�l��"� �Eď����_.��\��\��;�j���������EEaoG�~�Q�̏�Z����{ /��0h,h��s�nҎwuշ�x����n�:�L	H������<xӔQ�|���Kt���Ta�捘�3Gg��{�t����F�3="5�P��(�S��m�g+�e`��>�G(�,G+��Tu�g) �{^��u�r ��~ַ��^�G��:	���=?�}�Jfx8�,��ǣ8X���y�\��ugq1���1�8��,���(��h����b�
TK���+"���!B�jl[�g�(�y�6z*�-������ �51��b�������/?oߛg25�i0٥��ޑ��{�V@����v⽬lZ���R𔶀O�%��h#��=��
5̓�<r��^&�.��'�����d�k��TEM���4L{�4L������Y�L��9}MC__�������G�V�<=�%,��{�#�'�m�W��]�mȱe�G;������#i�9�KmՉ�.�E?j�/�ö(��AW~8�s���YSY7�^l�)���C|X"�S.82}��n����$I�� ��Z"y_;N�خP�9 ��F��,�D�p*]�'���j1����-�w�7.y�>�g2��Y0��c�7�0a�3'��V b�J��p�Q�-����#��=u�h�����+3յ�ZM$Y�|ؚ���i���l�#��RƝZcLŐu�{�"[�����c|8U:Y�}�Z�ǲ�m#��af��9s�`�i����t>���c�pNY�}x8ͱ�ypJ5|�[?�/��Ȱ����Gݵ��L�$�#MQ��K����$�t�184��؀� �Q��ؠ4�ol �<p��t��\d�j��O���,�Ϧ�����7��+���5T�S��i���QH2��C8������`���V���t��:"�N��6#���'&2BY��1d��s�bdt&F'`1�%öTޙ���o~fg��G�h��f���F3�S1I��ލ�3��3��m#��NB�#	�V�Z�D��iEo|ŋ��'Ձ��qa��=<��r�]�����zܳ�]s���5,�*�%�|���~�V]��<�9(Y+2���%�~��z���G.���͗�����js�Ե�/o�aY��z�JS+K��e�-��b�HF�L�Z���L��4�6`�i�e��H]L&&&2��P ���W�`˖-����BY&�SF�v�7�m��GN�U��ɿHw��-�?rZ�|�\$J�+���l|�R��ʎ�ߓ5+u��;u!sM����dHƈC���S���w���0Z�d/���+uÂ�p�s���?��q�k_��l�?�(�H<�g�"lG���HQ�ʴ�"-u�?�-��ҷ���hN����ƋO={_3 ����������ԓ���*Sd�:x�&��>�!�o�=��U+����T�?7����Q$g���ulذA��u���p"k%RXOI{� �	&b�;���F%-V{�5��F��9YT�[\�R�U�l��&
(Ǘ�F��GG讖q��'b�>��NI%sӘ��u�r�}k7"4�x��G㠥]�}�J���C0�~��M�tu�@X�^�`dlV}.���n�0���EG�u�dN��nY��}Q��¡�����4y|:����f����;�,{A0�����3R>܈����=q$f
�F���΀g��Y���� ���K��5�����؈���͛���)��ĉ�9�Z-1n�[F���#�0�ψ3��B{'p�,2�_�����(�Q����cd��̷�m$2����:��sj8�@\F
��m� =�2������Jӛ�Qd����֮]�9����~�D�i��NY n6`�6��^�m�*�8E�q�D�Yk��D����E#��j�5��n��O~�7�z�E�x�-�c܁��K0�}�+��*"�>��S�ч�S\lt֩���׮����J�ƶ�Y0��U��z�a'���o2TYL���Q����_~����x��%2�2%0�f�7�`ۂJ��,:�� �G�U	��V��K���J:����	)�
���Y���QTg��Lā/u��k���y�]8�o�}e=���F�x��8���U/�i�Z.�y)]膆uk�cxd�*��(Uo�'I5�*j�S)K��sv���Ƶ뚫W\Z�酳���ꫮ������3��e�:�;��;�,�e��<^�.- �	��sF�ף��oL�-�ok�i�ɺ�,uF,��p(X�e=dxxXzEh��>���~���t�6BF�c�!n�ޣ�c��#�&җ�c�P-`q�J�k�v��&"U��rl��N�i�d���XXSy:���eg�I��y_̶5����m��UR�
Lr�HI�u�	��-Ӑ隤�i�5��m���{�u��F7���rw�y�<�������y.y���8��б�|���+����0M�sgتIT]'�E�❌`n������^�Ϲ�W_y��?���	S�Ij�Ot��>,z�s�;�UC�_z�~�\���(���12����DnI&1PX	��*��L��V�υ_��Ȅ�\���k�D�kG,��$�vSH���"�1>��F����9"��!��B�����3�ECD@a���i�O������S`�	�1�*pD�I�\���2��*^�)\�B�nI� �.c���Jw=�(���|w&�K=7��4vf�흃��P�h��a�~�Ls�Ϥs�t�,�D^��#p�˞7m�o�bÚ��d�<,�ۋR� >�μ0@�R��񆏻��3��
¶����7�����ys���g�Vg���l�Ν�?�y���}��~�D����W]y�yCC��>V0!�v��Q�;&TO�����>��`�+�	H�K<(��KV�H� iЂa��?��`
&�+(����L(A楟}hO�IN��Q�h:r�4�hT"�{���$7�2���.�1>>���)y��1g�1J,���g��۠���Ȅ�%�1���������"*��P�p�X�)OR�FB�_�2▣q��ŝ�m�8�Ah;�����x_��m�j�u���>6+�)�Ϩ��Z�'/_�=̯X>����?j��k�V*��c�jHu��iP,�:H;�b���d���Ii>e_�����D3e�&T�.��ᮮ9s�%�j����c)�
�r����m.�C�f��
$2�ܐF`]Q�m
�ZT��Ob㝷�1�/��Z^�!�����,wɶl��p�^K"
�y��o��S�,,�3i���7���u�	0�h�0�����dd"F��E �ҲR3K�UN�	���Y�n�}��� ���t>�G<Fd��1<:��G���6üx|��WL�1��B�ulx�	�:��x��E�ǜZQ�_u�k���[�fp���D@�Z����E�@B �EIؑc�g��BO&`32嚪y2�ɋ��cX�'���V^s����G+�p��Xf�<�9��Je4�>��{B�����B�ɦ!\ ̈�A[���������Q�tEC���I�g��L���ϭ��ɶ@�����M.a��&�I�RK��Fzzz022"͉-_&�N[FF�h{��uns�^��hk퉋��6��`��a�&�����ֵX ��`6�$�k�'Biy��H$?<�|�?k��#���dJ�y4�-xw��r����9��Eu�Zg�~��O��n�R,�q�~���//Ɠ� jM�^)H���t��B3,��4����r�a{U��&�Q d 5�b&�2us�Q�J��F˃[(I*��5E��Z�F��R�    IDAT�nr_��fkX�'N�m�ꫮ=k``���
&�i.F&z����l���є�������
4ؐ��0��*��$1��X{�Q�t���EG�9&B6d��`r�M��w�'��nO�I~6:Y'�$�"KќF�����~alP���`�1jk֬O�o�B�OL
X�#L�dƏ����f�=}eHz�$Q����'B���#2���a�"�2�e�vA��I�Q�<�}��gj<�z�L:�];J)�Qa�^oNT�e�-ȋ�cl�?!F�m9OF�B)n��g=/{�3ex՜�*��W�^����T���-p�5Q
�6`F��P����1H�MϬ~�L�9�D���
�cc��]w}���_{Ҟ>�3��U+�9spp�c�L����A&��$W���8e��6)�H!C�D�U��g�aÁM�pߟD��t���9׵�3�H�5��7޵��O_�~O�I��Ϳ�fAi��A�!F"�6'�LXp�cK$����Α�ϦM�P�waxlbڻν������UAo:b��j	@{hO��	U\�D�*�N	��b���g>�¨��X�˺����<^����!��u%QW�$��;��m+�u�A]֛,����JZ�[���	��HPj9�
�yL��=:^��c�l~7Ҩ�j�.iΘY�7�[6a|d�s�06Ղ��(7�H�]���*B�,��,x2�,��IŒ�0�=%]�,�w���7o��㽧<�<�L];�ל188t�c�Ld=�����s���g"e�a��-�?Agt}�(��,
����9Y������B�Ê|Q��d���fP�$��L������^q��\�~�j0�nd�L�ɯ�hisz�7�ɺ�2a���bdhX�>Lq17^.�Gd�bd6���%=��v�GFǤ���\�1��⿙b�YAN�PdY�P�1�2!Q͘W���ʱ���Ъg<y?T]�B/{r6�{�=��oõL��K�
�@�Aj��g,>�)�S�h�����#�|�5ّT�HI��^�����X�3�UW9�$��&�ʖ"v&��Rۑ�j ;���\�6T��Raf�ݶ]�	 E���39x�����5�I��2�8E������q!a��	��6@R�ߢ*wˆm��b,m�F��ˉ1�.c��i&���}�2.�on���{��{�֞�ͬZu���QF�f�XڇB⡻V�e6��e~z��/��cl#d&�)c�Þ���q�	K���}ud�6����㽐�\.�V��z��"�C5�l�T�
�*�0m����R���u�����&F��6a����d��TMzF�����w�=�:='CXG��&W��u�NX��2#����K\W���%]R�a&*բ ��jc`hp��l�2���ˡ�Ӎ�[����eR��R���[��k�	&7����k�%(����Қ:��oA�����p����3p��:g�EX����g?# ���D��-Td���5���Q�U�Q���z��_���Q��9)�Q�x�́Yq�=#
EL��`:e�v�|�*��0[��b��^,�����.$�n�*�,G����̲4Fsr����8��@�Ta8.�H��L��1i��$(�cx�as��g�(�Q�ɩgt"M�a�(Œ6$�H�Ƽٔ�[�M�4�Xh/E�-8�7�v`٬K�۟�|&'r=)Y���'�x�E{�1����;ҿ�Sf䣤�x擗KZ��b�V�V��&׳a�,� �ı�#N�kˈh5�ZҬL����8S��v;J�����m]�v&�̅�&�P��sGjW�{w�g�7�Z$�I����(�(��D�����i��h��:��a�L\FP�����;�#`��س;ڈ�T�F��zhFp�=K�������m����ܦ�`¼^�+%Z`��j��\�yB�6���'UN"g�g��Lƕ��/��Ԅ�|�D���]bt��E����4%���Bn{� �D]0�C�L�>*F���˱�INQ4��,|�?��V�Ĳ���P��VLZ8���ba�E�[p���ޗ��(7{>��L$��O"8�S�����}���(B�۸����p�i��A�I���p�����g7�D�w�ߌ�~/�E�P���P�T�Nz���c��_E۪b�K��U49M�ra�1ʩ��_�R�� �y�*����b�D��F
�I(��ZF1X��Q	��8K�,�Fc݋��L[��E���o�x����%u�}EH$�4��D)��ߌ^#?��@��k�
!CB���`�'�x��v0Yq���ݼq��(j	Y�X@��f=բD��ObJ4��Z�\�#��ԤPK*���$���k��_n��I=Y͎אD�q�F 0�}�{���o�ֹmm�������%	��,��\]����c:):F�h��	��~�f��"f��L��gx���.���]�,-��L�Lx��hk�����v�)�w�X�d�Ty����jSM�M*��EuQdi^S�]01�J�矎>��q��^@�(�g]�;6O"���Āhr0��q�5��t�)
c�cP4U$Ʈe��U��d�"]�t4����8ѡY$��t�8!���M��=���t���
�t��x��BZ���f����E1�@� �ʕf��FF�-�w��1�8ҙo&wYXqᇱ��C�T�9���������
e�w#����uL<��>�/�+�]z�T"�3 7wF�����b��M�A�8�l��w�_^+<���֜�����
n�Ѭ6t���O|��q���w\q��oڴ�b�d~�K0����W}5\��6>�FҔ�y�5-�dJ@�o7��9&b{Q��}n���)��sN�����l|8��ŖܵdtJJ15
6#-����-X?�DT(�E�!�e_��"�!�(C396.�	u�8��ujlq�:=�z�K������S5*͢P}w���7���W�z�>�0@��0�p����e#4p�4R��¼�Y��+���6� ���0�)Q&������E��)�ЃB��k�\�zA��ܑF),-�a�(Gc��g=	'��碢5E>��[�����@}�vU��h��6���y-Y#�R5!0���{ZF~�p6"�`G?e���`��Q�o�60�;�̂�c��ĩ��;��	촍j4��s0[2OR\4�R��W�*��ҕ��c�)�y�5F&LA����y�BA�� �aH<��j��v�q��_��C��{g��k�8�y�u��,
eV�x��`x�vU��FR/Lu1�'����ɜjJggz��g��-�I�zl���cۈeۈfg��|}g�\3�":�|`
��`o��c�MI��m��F�S�OE��꙱��u���3.�R��F&;������KU?#��#348 �R��A����7S6�K���+��ԈlOWR*;�I>��� �Z8�����?=� X���:6$ݸ����B�"�T|LR�ʺ�Yˠ��bb��&j��0����Ŵ�NC����Vi�%`�h;]h�)���i��"�1
��P�`=�`�d�}�~8��Q3�p4���f]������M�a��BMoHm�Ѡ&�F;�0���/>a��P�k��&��s8�$
I �j�=��?�]�C#aMÀ_E`����6��8^����=� H^:�\	�S������8��3��vK>�&\K)0:�g�&TF=d��n�f�l�o<��?�7��|�ʫW�4п�f�HCT\OY�?
q����r�X@�	��	}���Z���a_��$ͻ{����k{��Do�(rC�_c���_s������=Ɲ���~~{@�+�U>"�)R�r�z*�e>� ��Ĕ0G���6a��F�g:q>�LF&W��뾳?�����	�k#��ER\j�L�b��%�0~��x�����#cb$�=Wz�|�=D_��f������I�zX^��Uo}6J���R4����U����
B�
G��B�d:#{J|��mԋ�(D�����N���]݊/�:K�u"P�:&c��G`$��"�m����bs[*Q;�0v?N:f^���p�!�d�y�wm��� ���Q�<��	X[��!򛰩� A�tJh�5D�a���X`�55����wa��(!@�5�6�Xv̫0�u!0+��nB�0S]������qO? O{���<#�@P*�g��\��Tp�?
����-�d�P��#�\b���}�������O>jWn�'�=W�������/RߌD[O�|A/U\��$
��ޞn�L8��(q˜ҭ�j����7�9������N���
�ǒn��w������FF+��b_�:�9Ȃ��T�]�6����p%� ����]`��-=��gg3
AıT�����ӕ[@w�)޶Z�t#_��ò��n��N����K�&	�����x*cw��5�����a8�o�v��}laSS�A��x����q�����d=}u����篗��\���|�� �jؿc�9-�dA'�,�1Bz摁r@0�a�hS���g��_� ��b�|҅�?��[�0fͅ�C1�N)L҃5A����
@��h�]�ܺt�[S��|�O`F#pӶ �gU��Y/ŘVCl�Uj��r�$R�V��㟎\��0_(�y�(�"�h��J�U x~��Y��F3�f�lJ, 3�|*>�I܎0�(�c�	'�����?���t���:><�Մ���N"�-<���AM&�R�%�	��������!ԅ�N�����9[۟�ӹn{��;�y����;3�;���>��k�Ѷ/�´"���W	�_�$E;1<ՄY*c��<�V��.����"�uF���{�%��zd�#0Qs��S���DLE���&y:�T��!b�A�BCD/4�gʈ���hewO�����7�>�^�f�-Z�'��n�}�B�[8=C��I8�̍&p��NơK��l����+׮�oX�T���/�b�&�]�i{�.-�^��02�0�#�C4I郃bP���T<���1��`�<f	ʅI$lh�{��}���u�+�����a
ɦ;a�(��R��/��!�Z��a,)!�+�&z�6���'���q��a�<�1iv��j2��4Z�I}��������9��Y<|:<׼!�P*��/�M�M�m�#�z����5i�F0�������VJ�?��~����~��ˮ����-�`��@����]8�Wҋ��;���e"����F�y}.
c~ EyC�yQ�Y6c�w֏��K�	�H�(9
�8�*�k���^��5c�����`��!�L�a���l!�
����c�4=#������m�X�!�	���~[:��)�5��"fn��-�}UӠag��b#�b�w�!�Q�gIC�8��B�\AWW�|��"/�N�02��n��whIt�a�'�q�����af��Cq�U?��Se�V��3?I0a���q�>��������(N����?���'�B;Tb�Q���R����L�PGlTT�E'�6B�>�����&nEo���U��1���L�����.�������v+�̍����Ī��e��b����.|:F]�z�j4����f�	��|���ÏE�ЇSq&�l1�0���=�i�j:�=z9�_�NE�����yM�"̔�U����Z�HZS9J�� ��'?y�7�Ew:���u!�l޼o�[w���a�ʕ׼l`��ۼgx?�^ �T��COwI�Kslw��J���L7M
�Ӏ���Q.V�1���m�+t�l�k�o������+��n_)����K�n��{���m#AӡЄ�ĴW�1��h��(V�ad�F1�H��i�U���x����B�SF�B���~�L�'�5��6�X���h �6���]�,�Ҙ��tctt��:�i,�z�|L��c,����#RZ����F�nel4���k��5��������ƪ5k�gǠ�1�a�
�����ߋ�1�AjBg���X5�p�.�}�a��Ui3�X�&4	�U$-S)�bs�-x��E���D�G�&�*~�.�E��#��"�Vo��?��Ǒ�U4C�Pu8F+i!�k��>^q��;����I�	�O����U,?�ժ����I(ޏf�0���/<
˫�戤�Xa����^5*��B��|.�(d�k��EU�ơ�:�w�k�ҁ��0��������{L��+W^����oJ/�D��B5�ļ���I�O؞�kh��\QPl.5*L���E���}K����7���� m=tՋ����v�G��F;H�Z�0���aK��X�WΥaKT;]Sb�t&#�/���9��ÌL&"�N�h&������p=����J';�,ٹL:(A��t���bdD�����TR S�����Hg��#
5X�p��/@o: �XO����_�'-DfuLRc�  _��D	R��9�Fģ�QД��C�@QfS�[u>���Ѷ�2D�o�Pv,�^m�	,��w����O���_~�h�2�Z7~q�(>�՟bE�u4��Fk��4�ؙ�^��Э�\�tLhe4� ǀ6�	�,��P/���k��~q�:i�)(�f�8�P�[x��Öt�Q4Ƿ(�eI�A q�а�ߑ��Zm�6�7%�g�OS~�u�Q��K:�F�n#c�Ӛe�N֯_�%���}�_�e���=���+W�r`p��
L�jГ��8F�࠯����'%<	`k	�*%�VD�~t�s��g'�ɣ1w����d3r�]�������(�/��	M�B�И��l:��]�#`��Q��ݢS�N�\5��?Q��I0�������_�B01u*��5[�~�L&6��p���^IC�h��}��x4"�G�Ea��7�Ӟ��"�1�?���G^p�F�ݦ�������q���K��|#60��q��⎍���-�E&!��I�K}I(A��f
�
�ka�c�a��J ��v���F$��6ˈzƈ/�
*1�&�[��Ґq�����y43E����=g��$ �)y�:~����O_��X��kFk��P�b�햤IT��@�R�X���; I��sI�?�ŵ��0�-�l�b����|�?8�����ӋFs~k��ux�I/�?�#�`4*�ʲ�wNÔȇi+i8ua����XP����９��{��KK �ß�����������o~ӛ_��3���~�+���8Mn�����$b-�:����뮢��h���MUg�u���i<6�_2V��~�2*�	k.L#��Ț�����d1�}%�(밣����KK5���Vh,�vRd��$Sg-��� OL���Ǆ<�K���ڭ�㱈�a�Zf�f�	&"��io��@QE��z��/IZ��m&X�t��X(��t��
��y=��h�R&�#y7m����4>z\�R�tkf� ��~����/}��B{
�Ě�/�f:"Ý�(#�����-+���)#5I�����MX�����EK�f���e6B�����4W�/L7���x`c?tʩ�1�fU�9,���$޿���s�&a��&-��u�����v���13jK텴]͟Ŀ��M�����Qꆧ�h�6"�í
���q�+�C�Ҡ��TqN|�G����IDz6)ڑ-�{�8�Cq��^����cS��,	$� 9~^�������K���-����'��#�8-��b;�'F&yW<�'&̺��N|�	}3u]��vW������C��=�qt3e�������kFGw� i��rI�����Nqֻ��Ϋ1�;.�k�o�:k/L��B[�ߝ���������c�7:�� T�2���Ps�������T�h���ęnI����S��y�Rt��K���\����>�ү�t��҄�A��1N��RaK�dys0z���;�[&"2���R�ϲ��Ck2�%G��z�~�%����Lf��η)�z���k�y�Y��몆?�AS+ ��"I�%�-"l6�DM���b,�S����K��W�R��k6$�� �ɦ��K�I�W��TR=    IDATf8u�$`���O~��ÛQ��ABJpl��\i���O����	�d
�Eh�@�
�&a[����qs=����i� �|�(���ab��k��ZH���2R@R�\.�J�H�$���H�:���絨���'11>% Ac?�exZ��j�.��Z
����ӆy�Isg���CQ�3��'��$��<�y�}��Z���h�L^{z�+W^�����k詊�<c�)e�U�5-F¦�(���kK$�ں��ے�#@���]�Q�}�oi z�벦,�o�s�{�����;[��]:���|��%8fR�0#qir��G��湶`u�A�-�o���(k-T� �چ��E&������ό�`�TLi�0�E��Q�/�en1�KŢ2,.�/5�y�P.��U�T込#��t��#+l�{$�2�?�K\�h���x�Cҕ?���JC `���H]�`��׼˖,B�ۨ�1~��ո�;_A�P���E�C�=�.���U«�y.��u=hn	7��v���5�t͑�m�-�#ؖ���%D���,�A�B�,��J΅��D ��G��ܞ�\@����V�H�D��o�15�^Vא�նl�R"�/r7�D	��k�
��ux����I/}�O�1���	II���I f@��^,���u�ѐtW����:��h�<<���G��:����V�k"ZUd��m��v�{���{�|ʶ��ʕ��cph�J��D&T�f���b2��)�ڙ)�J�b�K�����#�)I�))i�l����Ό������k]r�ȿ��?�0�E�Yҝ�pl_W�m��� ͛��S^[l��>i��	��fL�{���g]����,���@��Ta��m�(���ң���k&,�����;c��`�F�yc).em��k4R��W�M�qKB�|^G�9�Ӟy^�����4��[C���9�u�j��N#��(4�0�X�}F�D!i�k� E�ѡM�#�Ƒ��L�E��u�q�C�J�h����)�O��P�a�$(�A��b��%\�D2�.����2��͓i�>�(3+��0@��М�TM��"�k���;��8l��p�h��N:՘��$MGQ�	���vlUP�tz{
��$>���cio%+�F�4��j�,�jb���tJ����*��~γĈJ*jaG.kLt:���W�$����淿���ݰ��͘1C�����`��d=R:%0�$�ɦd��"M6��*r��z�����',�O�+m�wև�����-���}�vw}���mϓdr�s����%��qI����Y�����3��<yH����u?�����>?�6�2zVD��ѭ��Ԋ� Ɣ�pʕ���|� _.d��c|O���H��^0#�M(���k]���B�����P�����8��F�+6�;�6�����`W�	9K�M=,�s0�e�2*XXپK$����Afsd&g�#B�`Z6"��%3�"k@9�bS��6ô��$�F6���jB�r
�J�>�-$<V���1b����ɢĻ'��Ŵ��"FH�DɿN� ������Ϧ%�������5�J�(�ǖ�E���Wa�R��US ���t����S5��o�s�x�B5�8�T-X��,�c(�p�t���B���'A��4��[~��������AK�}���~��y�>�j��36o�|S\r]R�{Z>^��M7��mϑ�J����:����[V`:b�hD�U~5)�Ȇ�M�����8Ӝn;#��U7�Z;�S_'�ȄAaneS� HP6S��.4|7*ì+��X&a������Y�!2Z��J�X�J��M�4���B�u�D(ۺj��Kb�COQ�%OH)u����*͓�"J?�u��j�XH���")���e�\�0h����}[�J��2�j��ꂆ k�1/Dk���/F��2���D7(jz J�nq�!#�HzR�-3A�bd[���"A2D�L�e]�$��*��)�/�T7\��H�����I�ǫjr�7�]��gK�j� @�������i�@O2�1���$*eZs�Ș����d�1�G�2iϺ�z�S��U%�r��,�.�u)ͼ�-`��8n��W��;������y����'���_~�<1����������к3�	�C���������� [�p2{�;�x�똃���eQP&�y�d�Qb��T��J[Fǅ�&,[5����/�6e��X�����DD^%�g`���������ʪD�!�:U|Œ�L�(O])�Ƥk�P{S�#���u���G�f���t�ӻ7(/_*� *�-b�H(��$"�SdF����L6�������y��*@f:f.�'
n]�4bO�*��)�d�c�M���a����24��H�#s%b����<�����)*�p; 3v�e %�B�l��?w��Sފ�݀�E��\@�A��t�ƍ�<��>(�/[~ �,[��}P�WaS����ԖF�����ᖟ�?����JB�L�H����/:��~��f.���^CGD��L�tv�վv&����m|��~3&���������D޴(�#�	�6�l��s�K/�����1d�rMjS�&���d�RR��l�
��.���Q�tgi�Y+@@ꬁ�)�s�fS"���Ji����p,�h�[�#i(֯9���	Q+��Q��)�Y6�&G%R�0_��=��,H��qؖ��?�P�� f�&�R�UQ�9��L�vk�N�NY�������|�8Gm�ꖺ�����T�E�y'pY@'*S���7�i@J̳	�ѓe�9�1�!�"]��&���7vas�=�����Z���G��|Z�X��LM�COC,�7C��!l7t7�"L! <�nÑ��9�]�S5_�h��}k�`��~��!����]V	��[�s�-+�=_�����:����h�fk���A�ih�۽r�QNS�q���Ϯ,͎<��yٮ��_Ҭx��|.����R��~T�7{�D�,�l[*�����=��l�mT���o��]�|_�k;z�Ѿ��϶��%��M�l~;k����:�xz?�}T�-�׹}���T;��r[j<�֟�������3��������cF"���}y�mV$��VEW�!6=���*�	)-Z �K��00<4"�T���&�uv��u�&L�8���t�w�� HhU�E�0�8S9L�i$t~�F4�7����+yz�i�ҡ��K���J�^R`����+�'�����J�[&�N+�y��	�3 �ȸ K+T�e#����)%V�KDI�@쩨F(����91J�T�`��Ӻ�FZ"ْM*��&`g��"��-���g:j�p��f�Inl^�r�f�Bf�f���4@�v��R
�E8�E8�C����l�A��ڗ<IsT�f�6c݈���_���~��Ra�Ĩ� ~L� N�&�0���:��iÎZx������sW,��{fW`vv}fL���/*���$Ǽ�`B��:��+��Mcd�&�p��ehO��<x�R��TC�P�\�� <)���Q	A��fv���)T4�mc��BF�IZA��2(�@ќ��%{@,[�+ʋ�Na:��[bęBb��=z�|L��`NO7�'F���c�����b
��mUL& �ʎ!��fb��\8a[0X�����Ю5=R����&`)\ݔ�E�SO����)+�^�j
tKU��x&;����TM� T,���V�D�����bJt�TpE���r%�E�1.�5�Zo��2�f��Q.��_�j����C��D[/�,wI��5M�)��$	6����=nI��uŴ�#�U?��K����"��]��ؕ�0�ʏ\~υߞ�62!��Q&�֥C���]�"�椤yhi�4��lGj�|yH���&���)�b	�	��1ԫ5��"S͠��4����Y^k�t��vjbʋP��Q���X��j�cG)k"L9���4����#$fQ�?����#�}H��`�0}���
)�%�mZ��=�uކS�c�K���#Z,�U��L��� LҌ������[���&1�V���l�,�ԴB6O�����:Ua���K3�[P)��uj��!��F�D��X�a͌ͨd�q�(������Z�������d���؈ �S�"��i�@�[�vY�k��U6�S��ᘔ�!sNE&BI�8rY��?���v��}��
̮�������7�Y:���Ҵ�1-P#e
�����<LJmH\{J:ui,� ��Y��Ο���"w*}�;xU$'`0":���#{*z�j��ʸ����~���w��s?�u���yG?˖�o|�8��S�x�<T*�t� V^��#��� ]�"�A�m���o�)�^x�l�b�o���q���bd|�[��g}_����Ѓ[��i,֍�K���g���b~���Q.W����#���Կ	t0��j5�0������k�ӟ�
�X���v�������>�W\����=8�)O�;N�7,��?��O�~C�?<7˗.�i��;>�ů��_��PB�i�Q���G�I*��L�*��zX6�MjH<߽]U��mD�j(�{e�6����z�D�9� a��DA���y|Q*�?Cg���nK]W�=lS�&l�fr�/=�]�Ef�9��+�++0#`r�wn-�s嗚���E��=Z6��+�(�m)o�޻���kiMCO�4��(�~�h�S4�X�[�ItB�2��ԃ)������uXRdq��k�m�{^����C]����������kWI�޹�	_�������{^�/ƧV��5�����1�o��t�"�흧b���	�o����*��ן��>�7�t���/⧷��G/���}����/�>r�j��w��-�Dv�GF9�����8�����$�ñ/��z=^���X.���[�t>x�>|����m��|�z�4�Ѷ��%�"����W��z��8�����@���ڌÖ���>�\w��Xu�j���7�/�����x������z%��"�����;�2��Q�ߒ���,C�wU�g��i�IM��Qt���9FC����)�lx�ڢ�K-*F`������b��`X�����&`RTW�����gafz�㾯11!��U�1��(B ��ȪDA�(7�=�&�+�.(�1��=�U���ܚQ�D��<�����'A����ܦ�}�9�{��S���3$'&%���������.ߞ��&���@��ɪ�_^r��ɴg�D�:阃*p�zJ�����{�3p�7,5�i����)����GO����)�>D�����?$�jl���2Q���wݵ��U���K�ux���6~q�I����c��ȃ�đG�E���-gc���hۆ!���b�l�{=���sh�j�%,9u���0�D��؟᭷���G�sGMF}{7
����$����q�u���#PP"��(�Nb�XI����z՝X��j{�Ix왿㎥ˠh
Ə��0��9�O��_5�֥B��]hggXh�һ��(��X��n�Z�
-_)���tn����O:���oD��ܹsq���1�i�ᝏ>��$��#�'�����p
I騏�ըv�vZ�`�IAaX�����Q^�������A�_��n��8��}0����j��/z$c��utm�o�km�l�}�<1�����@���!�z���� ��~�����A�Ko~j����-n�_i~'p�@���ҵ�Ͼ5EbB���kJo��j���G6l�������>gҭ����eiK�ݐ}�+��t��Th���'1�f2�s@�c�>g<>��$,�=	�sv�� te��AOv���q��a���q�}ux����/c�O��{���Ϭ��@�����4(�v��N,�sث��p^�h|E�{YX��܀)�g��u�/��ZB�"��'eHoš{�ҹ�����0�O�QPV%z�T�ၻfᥗ���#���Y�㙿�%�O�xP�#�������B����V�ŋ��[��঺��qjf;6��c����/�)�:�q�4��屧b��x��Op��D�%Ю@V}�NH�A�N�p�D!S�m=]�$QCBp�f�,�H2ZZ.��mH�ۅ�emI�8��3������"�z����i��/^n���W^����RRY��I�A��8C	d_cJ��8dH�5�&������	0��#�'b2��O�3,I�)�l�\t���T��t�'�3m�qm����]�����]�����$BE�0�g�wm<�S�=bB���"X~��7f�k��Kwͺ
��%յ(.��'������Ƚ���c����nƁ��������x�����_�mwލ�^x���P�@�����ل����~�V���f`��-�EH�6
|���[���s�6��TŎ��ԟ�(�C��3�{�c&{�ML�n!�@�H��~�����}��~~n_v�z�Q�o�,U��9�L'�f!���r^X�ܾ��e���[�q��?ØKG�SN�ĉE������/�aG��F���#��·�:���#�V�s#k ZV�xG'�~���F���JKвm+ҙ��w��4����M�p��j1v�Y澵��[��1`� '�`;^#�]v�#�<��*A��)F��`ȵ��������Y�b�4�-L 7}"&�V��]r���AGZ>�@qHy�Ç��G�����S��%>�Z�P�����5��=��!1���Z�8(��UƟgށg^{_��.�{-��_P3`���a�Mu�6e2FChlh��kfA�B"�+���>�����9#f`C}��"@l���w4�cǨ��bݺ��˞��/G"K�BRϮ�3�݀�����h� �){J�#oE�B����?�^�SN?s��~��2'�r$���L���>�K�?�PI�"!mPW� 2�rB�[�x��%=�n�����lۊ��:�ɸ��+�Ǯ�0������Y7-��o�Cu�@̞3	�.�_njB0\�T�ꀜ~$&������-����"Z���Nq�5`� �#i��"2�(�� ���o�����2ۚw�F��|O�-~����+���j�ք���վ��c�C���}����36_����'�'br��oj����u%��B�f"������Қ���5aic[��C���{�o�v{vQ5v:����	���=�;�ڈk�<��� �B�.C0~��"��[F�W�1u�<�|���r���u`-�=�h<��۸an
*aK�!2�"���b��b�\s��@���W`�C�ᯫ���FH2p��s�l�������o��`ql-�x[3f��=���8�l{܉=�\�v�t$�ڱb�\�����櫸���`�/����J�Y��C�^��ڊZ6m����n�c&NŐ=��a�/�����짃0���}��1������-P]梅���ǟ��s��߲pm�}���?��_��"�݇�H1D�� �T�n�*�N�t�u��q��{K��Q��f�K.��ª��6L�d�e���i�[�-O�76�a�&���>ڙ������w"۵�G���v�І�O�Q���NMq^ߓ=�C�!A�"7C���0���ˣ�#�<Rؠ��ǚG���*b��������.���}������G�į�^x�>�:S�TDV&�x����wp�Y�Dxs�mO�x������0f�0�qX�-��T_ w�u6lj�,D[w
��\z�/�Ъ{�Es2YW���[���~UU5~ޅ(,.D8 cѢE���&Qqa��d&��!��?^t6�L?�7ݲ ]i��cGC���ґ��?��！�y��Z��Dgg;N=�XX�����=Z��P<��&႐8N+.(�B�θ�S!Q�T⍛�MAu�[[�`%:��g������ݑߍ3�X8����� u����gF���T�b�ecv�\<`��ճ�x,]�60a����/ۉ=����¢ɢ�zO    IDAT;���������Ϫaq�NU���ݰ=bbR�>��sM*��l1�C���]�(���DF�]<,�@��X�$]4!�3h!HdaO޺&ytI�dST�S�z�܅��,��3�p�d�We�����^��R�Z���dX���
�2a%O�g�m�Є�K<��fKO�x����1��)N��%# �m�4��*ߡibW�ѺE��26@�{Q;\�B�dMO����";���)j�H}3D >��b�.���(��ud����]���s���Y��ۙ���vv̈́�m�a_�����p��O����4hV�.X3��=��vv}�3��ū�ݝ��2�hy��>����؋�H*���@tr$�&�y@��$==�����XN�#	ٷ�Zۆާџ�rn��:����d�(i"�Le�G�Y�eLOQ�6E��,�%#+{*�4��d�Hg[+���E�H�;-*�4��N�)�D-JP�/7�9Ӽ5K�V�N�GCRD��0��d/9.���S����IC��`R�$�GD"��|4�32���X�NY����H8o�ֻ�����!����Ɋ�����wv�?ݣ���O�T��N�����w��U��0!;����=z�Kw���|�L`G蓇<ysMY�PW"kc���O��x��;����w�%�~�Kɴ�vT)�U���p�?{x�vZ�>)~�?Ec��mX6![��{��b���/Y�X_�ɹN��S3�$Q�4Ģ	y�VF]ҟ��=��
]�#�]��آ5�	���6��2�����S�M�N���U�N¤����Γ�&u{��E���#�"�{j�*|�,���%5���ig"a&d;���H�$�5ooiyy9ҙ�h�,Z��&**����l�"����d2-݊QGU(ӦM�o���W�����$P%!3��-|x��Q}�}�q���J�O�d�C�O�mY{�n�����Z>���}x�ͫ�w?�z����5V�ѣIQ����^��Q�-zM�8��f	�Hz��ez���nh�#&T���zlqd�1U���֒����������vd��-e���W��Y�!ckH��5�򋝎�C���,�0�)�:� ��Ue����Q�M����(UX�g��W�J��H$�&4#5ȒQ�>��@S�1;Ɨ$��A�2�9"�s�B!tlGnƙd�i
&̂��,�ԑ��v*P�l-т�����%�q|_;��f��ۜ�Z}�:`Ĭ���Ѯ�gt��]��=R�;�>������DL?�r�ԛW�&2�=�w�6��/��q�/�����稉v'��tHQ�����?��x�ң�WL�q�^S����AЊ#H�@�}�=W��/s�����t#T�4$MI�]
�#&:�"�+�&�)�OrC�j��N��LB@B
"a�7}H���q���B�f�P3�� ��W��5d6o�t���H�
�&��S�v���
J�Ȯ��&
�[|jLB�M�gVX鱗~1�E=K,rF�ݑ,�y�T"�u�m�PP̥��D�	�@ҋ���{aa�m�&�;=]B(�g�����C��q���x����DB��.�kɂ�L�I_B�wJ}"&��~���+���F]|�ڙ{����iuJ��R5�*�E�-�t�9^RD��_�	�w��)2a��"��(���N�Ў�@1Tl�3�B�KT�G�5�o�H�t�t*R�M��,+:"RA;���P������fNrqˇ���8ɩ���B��A�f�@5�t����d��Х R��tvII����b!��f!YGD��
�Q4�4���c(��dI]N��Ԃ2teT@	@��-�
K�@8 ����ۅH���^-�!(6����M����v��tJ��{��y�-�N�˿y�͸��ѵ�^B��z�1�d��󧰘�%t{�$�'b���u��.m��)L��W�1'����W��ˊ!��=��ډ%��M��ϴC�P�1񖞘H�L�DN�@�������ة1�U���*�BR��3�������(�t!$T8��,>�Q�ݢX�C	"-��$eP����X����+�4��>�(uY$�xRF����Q�T�;�������(^c���ƶ�Q�0��5�"^��3!�Y:)�!T��b�M��~?J�J�y�f�.���Ѩ؍�=�E/�lV|~���R�玎.C�3ݳf��9�N����k�{��.	G"�X��]��_�`2��%t{�$�'b�t���)7��I�?��A/8�˾�[y�2�̓\z)����S{B�W��F��VL��#��z���i� ��nԄ-D�8���|o����Hv(��Խ�y[	�T��`"����2BJ>�	�ӎ�v5���s�D���sL"3KY�����),#Z��n��OR �� ��x��t�'��d��.ji>a�&�m$Éِ�Ȣ!]�"�˲��3��Z�Mö���m6-9@��!7n��JB(^Bl����g��r&q��b�����>�%��w�Mїߍ_M]~�/��C F�N�������}9'��vF}&&W-�����.����^t��}	7z�8�~MS�S�#�Ɋ��@��Woorzx��X�+��	Y���	�}Va3�X�@�N@���#+���!�vT=oS����l�K�Bi��_#�;~T�D黆HO�H�H�_�ӡ]���d�v(�&Q|Bu���8b�4b�F���Ί�ӊDf[d�ы�2�D$�҃mY�aҜd�BBF;+j@�FV�&����7){�e���%h�d�qk�zv��,!��(R���nēq��K���\�.���ŉӨ>TVV
��BO��$&��E�+�;��}��8���k�����%%?�+�婅���/���;%�>�;�}�b�+7ӑ�IG�}����+�Ӗ��Y�P�	[�A1����[�~J��ń~ES�&ð�A�
[z��KiT�S��)���W5��idD���h.������('ؤXJO�n�u�$۞�eS+\�D7�2K)�d�N5.=�_4�,vU���4���4Ґ,	��#N$�P@���R���1ғ�E;!!@4�,;�f?ٽ'�#N8X�`�86khkC��aK� �hd$�=GE����j�;�ё�н��t�U=��s/"î�ȧ�a۳��;��}t�D��lքj�pؐ��O̿�����/$���蓿�w>�v��y˷d%��u��a��"���f]���M�P�¬h��,R5�s���w&$��V��*�vf�,�V�rUZ��O�3"5�L%��Y^^&
�(%�*���	���b�b*:T��r8I N��v������P�x��?(2�Z�nCA�X?��ũ/��`�Q�衯#�9��:�zt$qĻ��Cޠb�ެ6:���#6�#��fD5|aA�:��v$-l�#��pR�����.�_:3��#CG|eQ1�e2����rM��7�b�D�!GLD+]�SN:>0fL��ԦM�����5u�@��S8l��9k�]��}����i	􉘬z�咋��ߪ+d[7������z�/���r�/~�`��5��mK����ڙP�����nD�}OL*�n)i �r�5?����~�`��PЏ��� ���D<��� !1�%S/R���Sԅ��[&;p_�w�Y��K���7�������; �w	Kj�Ku'��´z�S����:g�(��e{�<�����ɨ��L)�@��c��� �������ARw�.�7^\�¾�ˢ��A�A�^����HP�C�'b̲�ra7C�W�E; W���NGn�/GLAbb$�{�w�K+���/��O\���>���GJ�>x����?�O*���xL&��
�>��k�_v��v]-B�l¯������_�h(������oxV
��c)�J���-��El�?�L�+&T��s��L�$b>!�[8�R�;c��v f;A���`����n�<�C��	5���qU�'uSdji�����վ��?&^1^|F��Ϯ}	7Ν'���Qe|��Ȁ"q��a��������g���9�dE<��ø��;D�zxR��\bıy��d�B5"��@��u��Gv�OO��/�n��x���#���V8����ۀ�I�d�������"��8v����8�h���w�����E#+ތ�g��'���Бv�_"<�H�}F���D��?���"��vv}"&w?�jᘅ�:�j?(zr�W\���I��Oˎ^}�]V�� a�"�ED%6�?�_�ߩ/��ױn���n:��V�WLj� ��z� kHf��1}�d�)�����q���E�Q�u�Bu��q���V�>���A�c�
[�`� ����͛�H�v&YaWB��t/��e^��"	EW{+��aÆ�,��"<��jܵ|�J��c&��Ѓ�Z%���%�i'ɀ�Nc��1BL�߇��f�uo���nX����vC}� �q�Y�I..D��]ɴ�8@�ѓ"��L�����7�]K�%1P�r��~ⳇ眰#��_0c�g��O4�Bq�G11�ލ�w��iM��	��b���^$&c��L�E�2iPo�dkr��sc��t�;�������Q�-uO:�Hfm񫟞��x�G�l���G]����;�zeIu�O�J�DX]M(
9���·��!�:c:쬁�m�3g^E� k۠v��+�I�U>M"B�%�La�}�����0��}��ױ`�|��F��~!>�8H���Vo��3�s�u�Yv֙�`��<��y�-��q�% '���(�˴�~#d��S;j4���Pte$�P�꾻���o�c,�i��3�V�@[֏�m�Ϩ':���)v\��)g���:�/&��a��#&��D��l V��Ɗi;$0>|ƢK�<�V�`��Y43�E=�+oZ3�Ť���;9�>�?.��3�C�dD4���om���sv�p�O��׻V�;yMCk�	�e%��=,ȗ�ҩ|H�_ǔ��s��ݢ���Lh7B�W�RL�*���)`�-�EՀA�~�5��$�����p���!k8G=��_@��P��`�W�p�U��vϽ�Ǥ)�ѝ�6�����(�'��hoE�PP{���#L��Hgp�ig�7Æa�c�GV?��+��e/ўĢT\E.���-�P�1�r��1n�~�O������ܻ�Y�D
�N�����t�jQ��z������k
,��O/gBvǁ�����v���T��2�����i8����N�����>��K��Ǻ:��
ŏ��Щ43� �ɐ���1���1_���>����#Sg-���P�'I�XPһ�e;'����M�xU�K2m�4yś�>�6��]Y	��Rq�O%�����Y��V�_�=�]ߝ���'���ùǝ�z�0)f�B?9��@a�Hw��EB7P�Ŵ�3A�;�~��ϙ=����	�Ȅ�G@�
j
�$�.��KQ���: c//���
�x�Q��V(��h����C`GGJ#�iQ�"ٺ�UdM��SN��g��I	cſ>� �^�~:*��5�xWR4��k>�	 !� M�CO&p��q�c��`�!!w,���kVc�AC��2���h��bA)�B[RG2�Byq!�]B!q�J$$N�rOeO|�_��H(��,��ŀս5����<rk^~]'��|�k��{_�*�eȁB�����	��\u���� |����L��ܾ��дE�%�V�?�l*%�@�*o�0v�я�9d��#�?3�=�t���Z�a�̄!C	D`�O�i	�����mE�2&U���2Q)�ae����Q�$`wo�Oʊi�����b�P���\��O�J<P��bZ� ����q�)	k(��I ��a��{��1��+��YaA/?�n�_5T#X��l q��j:	��w�����N������s��ڊ��"<�z5n_r'�Ű�(��ڭC����e(z'J��:�må�&��CGeT�~�����/")BW�BkFB��G�D�Mv-!�d�iP��B���ڷoUhI�àj�3=ފ���~|�o�O�l{F����ڿ���M[�:��`ka$-��W�FcFYG�Ja�%7?Yw������0��O�?uZ���5�.�A�&d���I壪q� ���8v+U^XU�L�^�3]tY�~�>}٩o������ytB���V�Z�ʾ ��hk�W����~��" O��4Ƣ�|V+��!�$`"(g�M'�����3D�/��b��x㍢�����ڬ��+=��(��P�t�8^:���0n�8詴8
{��W��E�j��h5��ԝ�4�����FE����F���q*�9�1�{�iܵ�> T���G��uYxoQfY�(V�(����#ٍ���p��Q)))��;��+o�#L&[���Jt�*��@�AM����o	�J:~˓��!Re�Y���T�R�͌X�=�|��"���j�ջ��iC���VE�l�<�~K���|��.2^���W@ĬHD��S|"������ħw`�A�ُ�:�����[� �}$&W�T�갂�e�8~�.��
�f�ْi���~U��#+�D�'��N�+�I8�R)
�R<$z��z~/�'1EΓc�Hc�}X6�(�,���,TW�`ʤ���(�n��9k�������@�;(�P�@��~#)݉���F_�S������Mu��V�N@�!M�&�P2�)�Q�(��?봓1���z����cɽ!r-��m����*��CGI b�ڒ
|�y���{�$	RA���y�����~k�FV) =��36�ϝ�C�%<����K����(t��|Y- ��&�N
�|������Y�Ћ�*�������p>�#@�;Q�2���43-vv��V}�C�^�߷��bL���1�c��uw%����$�:��x%t[��j� ���_�9��4��9�K�o��D��m$�}E ����-&��hF�7bE��ȴ�ѻQm���2��3�]E�����h㗘��9��*����3K����W$QSA��t�b'q�޻a�㑊w�������5so��/B'��[*t[��}�3�B�z��IaCo'�q��S0rة"v!�Kp���Q��~�b ��@<=�I�$#���x;��>�������ߞC��B��/Y������R�Oܐ����K��
[ٟ��P��DE����f�"��	�SR�x��3r�K����H�X�h����	��_O?�t�Sr��dփ�L�G`;�@��ɼ�?�Ϛ3+���CV��&	2[��~
�˚�*��e�zVd���!�$=Ew���7����T'��8���玆"�wQ�=x-����uB�Y&�6=�3���a�X�<K�xF�n�W=q�x�g$�nw~i��R�p�v�����gt�]�Qw�L$��**�����B���P�¦�v_:yuQ���ٴ��P5`vl�ؑg�7�#�=|��s�3�y�_ DE��CϤ�(���WW#�B*ٍ���0�ʋq��u�7d?�ߴ �=�
ԢJ�%?�R &�i��0����gi9�3��$s�|^�.��8)Ӓ$v��$0��,�C��ԫ�GlS�͈$
�Gf�BTț�
=M�0��ӏ��l�����WO����5L�	�{}"&3����-�@�Vd�K�$:�Ȋ�q���i�?������+2T��m�쭷0m۶$I�ezj�rkU�P�-5����#&��%�MIV
��)I�%��))��(�l�XY���k-fM� vYEś}����/��P���8�!�+#1U�!!(TSA6"�(�����X���7߾��/k�{l��A����Z0aYv�/Y%�����-����c�oOG2�K�d��m�C�F��X�uȧ�'�����m�UUT��c���������8�?FR7 �3f/��#v6�F���z�8G����]&�9�]@�Z�k@1��B��N̋�Y���aj�  
IDAT��v-b�# _��<6���/q�pHRz�\�^��W�uٯJ�6�l�����.���ۙ �y>�wN�$�ZJ�%����}~4KOvC-(�����k�r�����'���2W�Z�t��=��z��t�P|h��~��G_�� ��E'��!�w=����\���%��Q�E�_�����ԇ_�_�[���Я�?4Ɗ���7��~d���Һ_(�W�]�����e�G�(��Cc�gL�	�<��m�S��W���Cu�+�����Jq�ζm�uK�}����R}e��%�� ��jݴ�6[�O�B{�*�ˉ�]tv�g[_�Zv�i����GK�ԧm�s���~&���O��$�5j��8WSdzx?SQ= /������Y�y2d���]��磴4}q�	�|�������u���[���v1M���c��:��	0&�b��w����y�,���x��:vQ>������2�UsUe��������p4������XlC>c�7�,�m{���k��g��	0��� �I���yS���"���c55������iw۶GX\SS�N>c466^h�ʯ`[3�WW��������)p �Ȱ��Ī��:��	0&�b��w���Y9�o��UUU��0MMM����f]MMͣ�����y2���ɴ���O�:F|���yΆ��-Isc�1�g�"��	0�������mUVPa4WWUW�3Ncc�%6��Ön�Ū��3�W�M�)��W�7���qf�5e�f����i5n���(kZjԭ.Q"��!H͈P���Ӕ**�Li��TPa���(ԭ�I�h\ϛ|8�u������{������}�K��"��Zz��v͎MvO�������#̶��rr��Օ�S��eQr�yI-��L���F���^�GX��@ Xl���X�� �ʇ���m�3E��gn�!�F}Z;��x���>y#}}~��(�荨�3�
㈼9j�'�}�O@����,:S~��������� e�[�r���>����"	ȑ�?�����W��B�g�S+J�.��f�n�pg��ѷ]EE5iJ�fWM��3M��Ţ#��'��v��[��`����Qx2� 
@gp�������JҒ������:]�<z$D8�d�-���.�<\ʏ'���&����he!�C��ޠ
�Go6���/(��$���ݜz9�*�?�oEFG�U;<i8z]�N�H�y�F�AU�E�+5�����}Bv^UU�tx��bGEE�m�
ܱ'�WH}�$��I�0p�s�u0�L�9k��Г��4	1 SJ��?�8�T�^)�h���w'V��N7�{XŨ�=��-��S?W�&�!��Yc�i	t������d浬�hR_a�SN�???�F�� ��c����|� U�^Uu��P�\�ob�f���>z��� ��M�J�}����ؑ�[��n7�y�2��{
煞r.
���&UgB���L�&<>���-W�piB�*zg}}��!�3)����@m��%m(����B�e���v��>���O3�H*�����7�Do�-]l ���K���r��΀�ׯW�y�>/��_���\�B�t��X��ܷl�	Q`���A���s%Fh&�Z�oh{�����Z6����Q0 �!��W�-�HdeH����;U�G��\�Ҍn�4��z���*���W��A���E�^���rE?��yIO�lٽ�.���E#��v�6�|0�<��G�	?+FA��X__�����U�ePcY�G�]S�,��n;��)�s���|G�M��T �����oE"sjŗ�x؂C%�;k�s��ͱ�{|�ȹ&-0��s�����z-z/�M z��r�>#����pytM��~Ѽ��%���'�|���8 [�+pa������.B*T�Z��y7Uې�Ob�oQQ��}����&h	K���S:j�[ڲ�����!�D��7{Ejr����#,�;{�F����BQ(s̎�7 ��>r� �!������\�z�����Ñ8���s��E��Sڙ^��zzz��>~4i�$:��Ae�L_��DLVA�1�s�sE�a���u74���$�M:���!B�����N��]���-��7^F���Й�,��\�[b��k� )ĺ4h�$�l����fʹs@!��@�\/dţo���b�u"y4���Kc���jHZZZXC�P-X^@��9�a$i�����^�u=�']6\�"JJ�T���e5��S�F�PZ�k��q��
~Ā�Z��I�O�\)�����5�[�KH����Ж��(/���1����l��,��ar�:�z|�Z��+�7���=�*��;�I'�3	�E���f��س�=w�{�j�>��t=��)� ���H<'���%�_��3�����?����O)�]�K�N�d�W�s�u31��胿�b��a�$X���`�o���
�UuU-��䤺B��@���
ò����q��
��mv�mm�� [f��	��ͼ�pe��������TyS� @�\��4����g�i���V��S �)��Ti��.�оW�s+017��|�.�]p��v����۶�jLU�,U�����P.8�_PK   3)ZZR�yHS �Z /   images/cb4aaf6b-8f50-4b44-a327-f08934ea50d0.pngd�T\��6��-hpw�$���tpNp���$������:x���Oι�����Z�ڻ�����]�]U�ȏ��0P_����`(�˨�������b@F���}r�>P��u]a`>����M
�q����긩;Y�y��X�xzz��:ڹ��:[�;�Xg����yyQ�����>�AJ���9.�Y#=���+HE.�(㓶&S��� �NB'�4P1SM
�.��*�˗K9��c�������]?k��7}֪����D��^ �uon���U�ߟ��/�����r�.{� ��I��I-��sS�^��2�����u�V��ړN4-ٳL^W,��/Lf��}Ir�|��$7i´��l���Õ�g.S����MÞ˅{�����ވk��:d7W�kNcvN}c�;��g���E`������D����d&�x�~�#[��T!w�+��l�dR~������J�]~%�@+\���5��e��;�4��$��?
��"���/]��h���	a�Uo0�Z�B�������ě��K����F�]���Gn>��-�opXւ��b�ݏܩ~��+�m�'쀋��ƣ1$<�q�2yώ����ӈ��+u���櫏�nd�OE\)w���?���,5~�\iuݙU��\g�k8bX��w;P���of?���ҟ��¦ߔ"�����v�,`@2�B�X�L�-`)�a�!Ѩ�g��]�a����T\�(�j�	$�k�]��[��u�*�V�o�tSt"-�r|p�N�p;*����U�V�ޠ��d�a1T��8�"gS:	�D��z�մ?l��w���(�w���5�q�C��8�2�٧�����VRlQ�ClmT�����|Q@OX���;JY���󘙖��1��	�I�K�T��ש	8�C6���R�{���
��M�[�Pr�I���dyY!H��[���|�q�8;�ǡ8�� �5��^s�aC��$�R�hw2��pI"嵡���l���e�y�"�n[��QGs�1e}t;�R�	�*������a e�����c�pR9*qqr����<���lŭu���2 "ǜ59��0�H�N;Y�zH&yW�#̖Q��%3�z����J�K5�GY���A*�X��3%�ύ,C��[�h���m�Y�$6�\��`O&w+b"<�4�\FB��
p��`Nts"S-��a�Cy�{Q�S[
���u�����o^�Hz�ri�MҒ�Qx�4s9��*�a�N�Q\&��2�D�x��g�����؈~ą�Z��̚�I����
�����	5��"��g���K`���O�4�Waq�K�>��f��������ɨ�ά��.������!����G��(A	c� �j���	;�*�T� ���N)��h�cN<��P��*�9�-�x#L(�3e�k�C�+"��+���R�9��a�������y�̺9��{�t�4�3�l��@�(W�:��l8`�l[6dE�R��Y��ef�	�6u����Ye��N�_�j�g	-�;�7�N��~��� Q�� �rH�b��
�Ԥ>1'�OG�Db���E�H�Bڧ�pU*�e�j-�W	�je�I�K�-��X�u���cb.<��I��A2[��@{/�L�w�XQ8��d}�ka	����_�Hhj����U�R���M.vj��%ep��ڒ(�hAlwP(��P(��J]Ԣ����y�$��m���%��f)��*�%~Î�>���
�	.�~��*@�B�������+�3�C�&��SW.� �Cb<�}�〽��*5m$d�n�n&g h1�7L��qT��A3[��5�^�������&��]^�"t�Al�P��oPM-
Ւ/�R��#�!`���ט�k��������H�QB��e�(�~����kA'HRy�0�Խ1lЪ �z�4Y��'�p��cL)��S�@V�凝�]�6N�YAl�2>I��tY�{�V o�9A�0��(Ԟn�~}�%m����;}t�!ӶX")�C��᥌��sk�uU��(N0�w��j9�I�Dp@:�@��{��Yh��R��AV�0��UB��D^�B�)]^%���p�_Gd�b\s���,%��j~[�D
t֢I��y_��\ϟ+��(\O�wǻ'�u���fx9���2�����oe}�Z9ff�A���Kp<��l���qq4
�E?@V D��{��f�ÔL�a^ht%�k�֊���ã�nM���|]�1��}n)�&K���Й��c_�S���f���!�ML����gy(�De�Lvöb�l����7y�ГSU���LV���[��G�2�Cc��`0�7ŢU<��^�k�����G�z+w����*�F&�'�AL�'�T,��Ğ���|���LOG�x�ȫ�+c
>}'Ք�@3��lo����e����`pA�t��q�7�f�D1�������~�������
'8�>_[G$j�#0�|�0�gJC��pd��� �u�yCт,-�/��c�e�L��$0����0
�ᱶ��>]�¹rtR9b���+�D���T& 8�M�2T#?�Ӱ	P���)��ϓH���Gհ�zzl��Q}�bH۱�û��Os@
�p
r�x������o2�wBɒ#ʨ�[jM��8 (��Q�oR�(�Iiuyy��֩�{�b�xļ2z��K��t��c����uؿY(kq��}��;�Bw��9���.�#�e$���85�~��P4n��(���3��y�M���NYG~@6.R�7:"��c� e����+^ҟ�BU�����0pc �c�o��;-�H��M�4�e�i"��R��W�ӫ���~g�h}J?R�ӏ��S�Br�ݷB������@����z�\�ʐ�9�e�>���&ō�Vb��wv��{ �*��	�%`d AW�q�v������Ծ��&#0ǌ_���E������<��*�ޞ� �(!CO�F�x�"Rn
�i�+�5�1{��uK����A��к������n}E��|��a��R��XA���Ȁϫ����u��e�$�u����{�f�b��j��L�F��
��vN�>��y����t7��U��`�����>Y��ף5K����,��w����oH�����_�[�����;�{|�ȍ���M^���UW�|4����� �>��h�.���?����e�B3l�+�Ӷi<f(��4!Q�^{$Y���Y��k���V~O��`��z|!�Eh���P��0Q�T���lvCw��/e럜Ϛ��h*a�G� �d���4wM%M�)������=����-ɌL�L�Cd�f�X�M!b�O+�����-�^�ҫ

?i�jҁj����eS�k�2��դ(w��x�s�$���&��8.G������o�%tޓΟdG��1��ءq�C���]�6;\���}c�ǉ��Yc�yoS�g
��n!1ywf ѻ��$e��<ڌ���zsٟbOi���y�wU�F�[1h+.m�Z����[֥~?%r_���.���wb&Y`�n��i�숹ƣlH�@K��#��q��j���* 3�˼��c0r�z6hzp�~B�9EvSP��ȍ�v��c�ͯOV$p� ���*X���j��簤�$3`�$����E(T�A!�o��b�5��hYd�-n��o�Rx���>s��?�1�ne��]
T�� xL\��d/�g��ߴY����W�t+m�>2��A�l��I䆼���ۘ#��bv+�)��h��c�������5������8.�:ű�g�١�ɀ�&s�4[��S"���-�2��(�p�-_�&|WR쭂t}@�}�I��o|�Z"��Ee��U�� ~��;���f��ƒ�ڤy��
�_L@;�Ex7o_M9Y��1�����f8��F.Ӻ��[G��VfH.�@��������{��S4#�Nz�O[�Ӛ&�wi�����cJ�E:�!��Ev�)N�����Z)������U`/��uǟ�z�!'<�p[��Պ�^��헇��'��2��(��S�ws�͛����xw�9��J��md>�l��>������S}�d@ײYa�";�2�r����n�MܾD^�т[!�x�μǿ�ݧ�����ȗ��{����hܫ-��g����̪�H:�Mya��� ��V��4��D�CKf�ꡠ���Ţ"��]d�������R=��4<e���8I�����I����*mc�g6�]΋���;��5����^j)T�x�؀�*��Q���,:�l|�-*,#ݗW�*�v�;<�7��x���C`Vͻ�[3�S���/�fӣ��J��Z�o����*�%�9O�ߖ�,J�5N ��F�KwCn������9���~��e��B��5�m���#��Z�x��/�$��4W+�l��o��x��2Ɖ��
<L�n�"d<��X�R��դ5�W�d=>k������*XŌ�6��C|c��]�/X�����\#��,?�`�$؜�s2�)���h���3��֯�(j1�
\}K��eUh2MGך��o;�@�Pܯ�����l޽�m�r��w��2�i@YC'%����g������$g�N�m�c|V�z����=%�N��tI����1����ʒ8�fw3���W��0Ù��ޜ�=���I.�I�54���g��4Q�\a<V؂s����[-�z[�e��9(�X����Z�*a�X�r�p�R	~l?�e9V�����:���o�/wx_xUЧ7���r)���gU�W/J^��?��n�E���7�S��U�Qz�; e��	����v�����y�x����N/Y�F����Σ|����&5JW�o�9Mr�)_,�S�kU�0�C��R���_S�t�6j�t���2�K�v���|�G�J��e�|��9޻fx���
��4Tָ�E�W�%�����-F4�/e�	G�蔊=OFr瓀��BܖQ�Ĝ�~(��i��)�#VZ�VR�Rt��b���it;Y3�A�#��z�Ъr�6�<@dN�x+kϹ�Ad'��_��h�U�-��U��[ E�y^*���k��-X���>cpAA��
�]~��y��T������:}��od�S�~"��,������Utmx-�i%��K���L�4�F�%a�R��Sʔ���붝��̖�c �֙����H����W��v=�+����0CK��d��{�b�bЁ�%�ѵȲ-ށ�K����.8���=%�sM�+59 �
�P]�$~�˲���O��=޸�u�r�*��_ݫ������\j�]���r��N��)<����=ޞ2��xK�s�\��q���jC}�n�R ��7�	aת#�<�`%�ϴ���(7OD#ބR�%qN�-�ԫrB8��g����Nk3�����2m,�^1�?������� �<0r�Bq;��K�
:�`�$/�!��oQ�?��8��򞃂��MOLP�(׏�����MÊ���5ߞ�~`�$���~�[گInUE�%D��{�Yr~�2�������ਐ,�z������RVr�/M{p;(�`�0C5�������R�4y�g�������\Q��G��z0yJ?^�Ni|��E{S���R���QWl�I��fK�Ę��>0�� L�����@����3���Ih.�-�V��e|��"����߄�_(+��2�ߓ(i%P�ӵm���k���\��u�R+.����8�4�z��M����P+
D��t�ԢYʹ��"��}ЁjQh�JkXl���J}i�喘-8��g�P�I�>�zU�M-G?��L@V���������u�5���[Л���Е52Z�U��U��"��[1'�Z�\��d}���es�Cͩ�1C1�F�/K�x��ot�l[UE���#P)�y�g��v�B��nG2%�ݯb����!�	u�6���� %���tc�{��8��V:[jQc�I�`�K��� �K-����_����,�,��Y���w�wL.n��C�� 1��A�s�ao�Z~ڼT|�y79A|1�T(�D*-�劆Lв�{��u��Jp]�������,�H�O4*�:+[Lu�q�
^��t�+�`��,T3h`F\JAa2Q��=��w@��Pw~�����Xn�����\Mm��w�ߋ��w���ܝ��1���؛y,7פd���dSw� ���9���KU�����ߥ��B-�D]��Y��$��+r��%6�4��}i6������Yl3��e�e'%(�9(hB�ɽ��&z@�#DU���6i����&����u	�1��X�{8��\��ڼZ�e�_�jf�#@և	�:PBF-�7]��-'��SK���Jݙ"C��-��n�(�Y�D]��|hn��zb��w�cM���m��'F���P�fp�4����L?��7F�EQ݀W��V^����S�J8����?{��;����o���3j�;��O������e�/41�I�I����w����xU2��ǯ(�{u&n/�������F͎���sՆ��9�����Y���z5��WC-�j�<��0^Y�o�&���,!6o�R���7��K#,���)�Z?�2i-�S��= �L�rǼ�ѓ�Q�ZC:�]��I%��%��J�M�������Ľ��,�>�aq{C�ɹ��3����!��*�����{��4Vݤ_�_���������bHp��d���x��"�xZ0�3��;"z')�,�a\�N*�Hǒ�e�i��`�kE�]�]Ø�*[�Sl�ª��gU%2F���(o5h\�b���x�)h�,�fG*��!qu�y���OL$6�9�������3���d�A��>�I��*/�j_g>�S=Uq���~F?�B.�����1�.�g~TU�˹�}���'q�5.��$�Mm'�)D}Y�ć��4��v��o�&^��� �Ӛ��7�R6䋑4�����]�����b�YL2̟ӳE�������t?C�FR���#��=��ݭ�ug��:yg��Uj8�ihh�-ux�6��W�;S:4-��ca~��\6��MRk*e��)z]�������#���C�)��p�S2����/]��eL��l�Zw���<lT���l�gi���s�hW�?B���5��_�|�,��1^�&H� *,79�($���/r;���-��c@�n�Wh��ܰ�ջ�8�i�)��BӍ����+e����J��%}󷔟�٠i��s`����7���:�o��,��U�JL��Ѯ��'�U���x�=ɬo�)mT����4}:2�]�-��ck50_Zi�Ӯa�� e��^s���hs���7R��@���{��mʿ:Di�3�J���To;4����-�h����kY��χ,���8?�-7��8��n�/n�۵P\ ��\����a�,����{V�ÁI���";?ױ��ї�	fAE/�k-3�4YNH6�|���
�F�.V�=�j���z>��>`�}$�r
��]4	x���n���G��څݯ°�c�u�o�C���؅����(�=|��nOEX `9��Iv��hD�Y�u�u]�d"ʽ{��_�,��B��1��lA���8O����V���֎�~{�5�A¡�|H�����r���P`7���vw�`܁$|g���^���d��n|�)�o�5����Z[��5�?�G(��W�n��=s)��sp�eT�2Fn�%���i���ŋ����w��	�e��\d�����v�<�!� 6���d�i?�t��s�o���f9�Ic��<,�C��Y�\C�w9�)&�-�����ۣ=X�&%�ȧ��������A��I���I��d0Zt�74aN�~��ɕ$�>����5�8�X��=��y�YO{8n�!��S��`�?:/Z�v`��! �T���/ ���m��A�ma��vP*�e�xv�p5�k0���kW�7�/l`����E�i�Le����X7K��'��ğTv�~W�=.�`
Ƀ�R�v5�"[�X�����IP4�g������Mw����]��ͪg�Cd?u��HA8��7%g� �A�?'پ�>|�:�ǂi���3��q
?�^È]�Q�����zى#��%��)z��/��dخg��O���ah^qQ�C��YqW=>C7����ҁ��cv�����E�)�9�_&���y?�قy���΂;�O�y�ar��8ޡ���&���e���=nb �P>����1,�Ã{�n�k0V�ĉA/�;c,5���Eqcb��gO}h��@���5��� ���V��~xAAX�ŀ�Jn��ة?��r�h�R�S���H<��D�1,��y��+�Cs�F�?Pxm}4��<��#j��zQ��]��`$3�T��R���:�wY�<���CS��nl�)Y��l��9�;OV���C��Q�%RM\��PW�޻?(�s�x�=[�:�~�xY^���<:�����n�~��CyOf�R�����9ʐwy`����Y��#���J��\��k�"����C��c����^�������N[��n}��$Z�v\�{�^�V*���ۢ|ѹ{r��ӠW�Ƞ]#��?%��z�;Bl�<��+M��v�[{���-�Z���_��n0��]?���s|i�[>i���e?�"�� ���V����y4L���kt��Ô�:�%����=5��ǨK���E�+C�������ԁa-Ӕvu5o|�T��?6�VQ�4����Yc����w&�~ga�fހDµ2Le�N���7 H��ز���q�&���7�A��������j~���wC��{;��{/���$�"�!Ǯ�3���S����˲C�w�IB8�9>�4�����\6Q��������$�ذ,��g��������
*��V��v��UM����ݸ��rM��o2�χu��ǈ���L�[˭�aV9��\�����с]��4=���-fs,���c�e�r�_e��d�p�d�MAQ�o\,�%h	��)M=���.��]DnL��7D�`���Ѕ@'��gY��G H�#%�	������?r܍��s%+4 ^�K��"�#���r��m^�U�:�/D6/G�}�0bV�r9Z6^�3���3��"��8l�F���}Z�!~@�_�����Ó9����`����l6w_o�2�2�{�ָ����b�c��#�km�������T�`⒱^�a��Q��ƫ\v �k��Mj756�׀j���o����Q��9L}�<t�� �[��U��7�i��w%{5V˪)�e9�|�8Ȍj׏�RT )�y9!l5�'���RB�0�i��DA_�C��P�Q�X��D��p�a�E0[@ě^�8	��צ)o�9�8���$���򚾢ȼ|���E�o�9�XO%�Cq(�[��#��8��,DI'9����#�qF��DĜQ��^�� ��	"v�k��A���4|mH����cM�/�j��{�`�D:ך\
v�|�L����	]��6��	q2~���:'���l_�f�,�@_�{���hL�U-`-.��w�yY���@��A�^�tv�^/��b���݆t���C�R�R�$4�a�D�ߩ"�ϏM�w�$;ju�?tB�XDw� �B�ݳÆD��m�̰d�8���֘g���(��R��;�{����8�'���}S���4o	�J��y`F) >���0}��w^@�n1GJ� ��A�gnCTE�w��z��Ik��0
���:5�0kL�E��
zHWꨩ*���0e@��|��A��������~wF�ܦ��.Q��hqm��!#(٦�2ל��=cɤl�d�6�qE�9��Km#�	���Zz�/������W���'��T������G8�_*9l�~y�N=!ȍ�	��q�=|KA&��	�N��U3�m;�Pmr	���s�Z��O�	���A�&ޔ=�i�$��A,a�\�=0Xܵ	�)�h�a'6�汵'�B]��`��4�F�(ߟ<����y���؆Ɨ��x���bi�D�j4U6�}��z����C_I�[��*�X�7�Ħ�=.�z9ξ۬Z7SqdW�5���K'n,g��D�l�����W1(2�_^���5����VLS�b��H�����a��BpD��۱�+.�����]Ѧ�c��YE��ki���"�[�������R�cbK�� QQ����pY�9�{UG4�L��'\������s��s$M߅�����Ԑ���P���Ē�Љ�#�o�0�6�){��[�f�5�x�Po���� �����P�V=׏>�0��ب�^i�`\Jy��\�Ee",[Ʀj���|�n.�Ve����KK�Ƴ�ȳd�U&V�y���i)�̡��^:�RςEoE��t'�Z�� ��!�{�Yn/��C��e���3���q1X�Δ���`�/4U?n��i�\��_V�����0#��qp�ngF���p�pΔ��ά��n�1r܄;3�C�k�m�©�hԳ������r>���P�,RE�z�f��]#nK���������x<��Ʌ%!_1�g��J�(�߫�&��/%�~M��|f������:wO�ԩ�e(�fOq��%^5�UK��ǂ2hpI������E��J�K�q�9k�5)Ͱ�bW����Q2�0B"�\{��#��Z�X�q(C\vb�a;f�`��ۣ����.��!V��*B�h�����6B�z�Cݨ�C<B��<���k ?�TN�n���!��&y�MnhN;�2�R��v�����BQ�r���;�yv�I^��{�N/�cdJ���!���5���ޖ|�v>t�O&�mL3�Z
T�8�̢~��A�����R!��uhT����w�1,�Oz�`E)��_K��!�ERW�݂a���z��D��E�����B��s�΄�Ÿ'��5=�s�y҈m�:[:L3��1�Uߤ{�j`�"�v��� ��D�|����������~�Б��碗3Ӿ!�z���3���f�.��}�`u������!����]� �B��OY�m��o(B6��^���8��N��ۓ:�S��bY����{l���X���E�Q�����ˈ�`6��0j����W=���N��7w��S[b ,� �9Ĭ����aG�E�TtKQN�(`��Q:����}z�:��ֹО�����S��3��ye�{B��-�"���$�(n7�F�Dĳ�r��ED�]��g��vW����ˣ0�J �.�}�I��Mts5*g�<�/,~e�F<ܴ�P��k��]�9�uH�?D^X�}@��fD8�t�H��e4w!�/��L�~��}�Ü,c5��8��������T���T�}�p&=���,�(k>o�`�(�I�1	�,��F�a�j�֣�i���!�G��y◍�'T�&�7��f��.F&d
*�-P�m�W��G���pyg���`@ǹ�d�d���}�.D�^��]�R���� ��!��:s�����Din+hQ@`�E¥@��l�!S�=qv� ��3e:1�?�V�N7����%�x�4����!DN,D��NVQ'��J��0alW`ݫtu�?Ί�I���xRq����*}
%4,C�����w+�{P�
�h�\������#�{>2���L���㜴�_lz�ݣu�]ѕf.�y\7�Q������t���j��F�F�YbHp~Et�brC��<l��sU
r�����kؔ��'�6*H��ɚ����먳<���gG��+�$�	�ͳ�B��O�8��A���=��_m����g����|����bDR�W�])Ym�L��Ƨ1�Ro2U/;O�j�*/���?��b;J
o��Rqe�/$��;�)�`%'��ĩ�z�K�z��ᯊ>��!!�#8ûm��g�]���/�/�l�I(j݆[��r~ٲ��p�%�#Vء�n�i�v�.�E������1���ȹ�[gd-J��O�7�HV�'��,2�@���>At�V�*iW��8�p����)�\��A�?/6��p��P|�`�D��&EZ)�麁e��m��Ƶ�����q�`���a�,�M�������Ð;��,#�<���MU��#Ƒ��^IL@g!�rp���1x�h6������4�0��r���w,�Z	��1��KYF�h��{
*�@����'��a1�M �g�0U��8������{"@�Xa��:F��ծ�Ӗo}<��7Xk{C��y���&� �����>�Ĥ���B�3�����0^�lf�8�[��d��jXEC8V���'��x`��M�Eo�}����{(�Y�%�uA�� m���~�n��I7P��H�x�u��4{�+8x�Hp`�E\�N�:IQO�WS��h:?���	A�p�M'���ߝ(d����e<�B�o��B�S��|28���'=�/6�4'QA��H �W�4��Pd��R{�{x͆��1J��8A�t�3	�ƌ��V�z�ʄ������ozt 962�<f.gD9�yh�>�`����	�z��z/�K��d�Pzȱ�3��M˔+�|�j5��(Ye��$��	�+��Z�@���*�K0;��LfZ���� ݼAfj�]�aH����@�7��g����֑�b/�$������t0z��T�ImP��9)��-�l�QMe��l�[����Qt�GՖI��ע ��;�������)���s�X��fN�V ~?t/#�h���	$�y���@�0>��62y�6�-P�iqZnB��L�Q����EO��NG��d*��zRzȢ�_? ��Jv3�ʀ{��HZ���#�%�V\D���a��]��~�5�3 �+BXfƎ�_�{�29�����84_���nm�~>�x\��L��,y��$:�N�"R�;+$Bp�lF;r�l�a/� $`rNJ���8�k��ih�ksb8��x�����Ė_V.���wc��(>]Jˀ��g4�Y�|p��,��|�S�k�j9WX�K�dL#�&7����ȸ�o��C�0ɟs�p�^!P� �w	�4��[�a�|&�uDDM� �ٌJPKȠ��A\#t��ď�|S"X�?��Q��?&Y�8q��b�F3�g�i�hu6./	��o�D�m,���<�RR�D��;���ȿ����� p��{e���9r7�s����g������F/�6)�Ӿ�~=� @�ix�J5N�a�Ċ}�u�q]�3�-��#��@u��x�
�ǽ�<���wF��K^<�M�Z�Q�/��[#���\��C�����H�ϒ��c&y#采#��h���vAvC;6Z�����z�x� _W[�Yk�)B6e�:�{�჌"�y�d���{����<�Gd1�m�*�Fj(���C$�2p�Q'� ����"5�r���'�MR�y؃�O�I��:�S��1��(�0� '��?�G{���X8��>�C5G<Q&��N���9Q2���'���q�}���U8oM
��8҈a���:K�]�����5 �}�cQ�z/C��0=q��zZߒ�6�u�~�����g��(�-N�q-���<)�����nd�ǧ�W1�MK����yY���B�����}���ٴ
�9h�@�w�ش���@���K�Eǂ��lJ��߿½;cݹ]�n;�n|%��'"5 �e�ɑ�H��Ggȱ�c��%��7��٧����`�,��W!��Eg��c�	O��Q���5ǥd���[I��@�	��k�=Ba�*�^�����P �u�$v��Fi�;�Y�Z�*�LWkf8L�y����t{�ܢ�\8�7�{�J�[�O�-}�=��If v�,]�9�����X�{�HW���6�<%
>O�2	�9Vj޳�VƖ\]����Y��.o��qy��}�#F�����s�%H��,����^}F�""�p�X[��U�}�p�2h���:�v�G�&#>���B��8��Q$]9�O�d�vs�����E#�=QXb��T��@�Լ�52��}�G��Ȫ�C���xH���3�]���@�D�\�z������St��=U+)��N��7谻s�=6Q�c�W�ȟ�.h�R��ᢞ8_�&�/���[��\�p0/$ܒ`S������+1$A��dd�I�H�X�����R�A�P�ރ�ѳ��a/~FiR�M$b��]zV�K��3��3��y��=�Z�f�	�yo��9�Ft@b�������[ R�Vg%���VR����vKk|��ss�z?�Q�����S=��,�u�ӴI��w��-�,גz�)L��n�������;�Ѫl�^���&���֎���Y蚾LYW��!�X���C�^������^� }r�yzn�z��N�+��]�a����&j�����	����O����
_쫦����
���xen�hv6Ց� ��L���Y=�~�s�Nca����!J���)>Z@-@�/^o�eXN�����I'�P5�R�%�z�'o��1��}y���"9� hF��j��qv6�J}���Iӆ��/I;C�K�-~X�B�p^
#����5A=�N�p1p?\_�jDj�d�Es���Z��BԄ��v�l?Yx8�Rd�ۿ��f.'I*ӷ�U� @��`�5�� לD�[jAj �2�}(����`纤x����kd��`3d��r�é<Ck�BTkuzX�Ab��`�Fl�+"=)��_Tt��ǄY��?�����/of������.Ѹ�D��E>��-�o���&2O���ۯ+�� nL��.���dO)�ش���(���7�B>�gs)\�֦���r�R:��L�X�g�-r�~&gL���[������� ȋ���4�	�e�Fo�î鲢�k
���.�EǦH���b%*����*��P�����������[}G;Ҵ�b����#l�ǹL�
[�5K�>��c������՜��h�9��˯l��~��|KB&歒@�Jgo��kpr��K�C��U���L�ێ���/�GLmS3z�j�c!�2��;��|ꊤ���XvgeϦ	�ˡ[g��.o�1vJ,X2�\���4b�����#��8|��ҖP_q)�
P��FΆz[\[��1�G� oz����;��	���]��'D�@-�ET8�-��H�S�螞$���wB#d�&�'2c�	�?3�?������Ի0 ��v/ۼ�Ht�%9N�$^��؇��z�o�(�PxKNq��ao?�gVqyjŪF��d�4W�"d���wCF�h�%$�_�)����nV��4�v���O�<N�s���5���O�=�;��(ReE���?������_ F?`t�8'`��E�@9�L�	.� ������6H����&&�T�l����:�`\�,w�a<�in>FG��O ��s�d8q�X;��t��M���4F��'��`�b:�}�N�،�C�����Ww;qg��;@�}|cО�q���<��C��4�7 �l�K���S�Q����ʒ�෪=�^�ڰ;�%C�`Ze�_'4BN��bK1�^[��g�[�ޖ���c�k�7n���/aT���z��`[�D��a��*��z*��+�ZZ�t4e�������`+�W)�ȴ�ux�d���1t�]�����:S�j�A�J�%o�o�����y��݄�7��R��GH!`�%�V��G�x;�ɦ�
l1d�otN2
b����N�pk���I�f��v64Ȏ�K\��U���Ρ���#�T�ܲj�V�X��\a����][Uyb�:.��MM.�z��:G���]��A��y�
Q�ů2��+�x�
�O�f8���ROJ+���$f���{��T=�����|802uN�G�*�w{~V�ܛ#s�����;�{�:��:+b��4��VQ�a�q<C�����)+���CC���8��iJ���ҁ�y{���)\� ���8��_�$3�����cb'�=��dDf{"f�v�8�u�&�OHq�ڝ-n�%5�E�'�AL���_�B6LD���U�(g�7���M��^Z��Rco��H��Y�3��c��?����ϊ���ꑒh�H{���˿A!{��I��(В��ͶG�1�^4;�a`~C���_�M9z��Z���)�f�N@:�pg՝��.4�p��C'7���Bz��ʫU�r�����%�
[�}v��P�m�� ov,%����ىQM+����DT�K}�F�����b8
�t3��x�{�t2���`���GQ9}��9)6�c�0���a,���=�ч��\��$	(�*,���K����T�����퇦?Lڥ��|����i�I�}z��ȄeT`�c���G@��x�@��t��Ş�Wh
h�"<Q
���r"���$M���\�ld����*�����2�-��k)��l��9�C%)G,�yҖ_����h�#�\|[�3Q�[`&����
��$0Z�q��{6*�!�&fpk����^���N��-�ASM�F���o��P@`� �ٖ"��TS���k)�{>�q�%��B�>� ��</H�Tw/��z��t����ǝ������[���))���a��KBi)��n��.�����Krh$�~�s��>��'׵�U����뾷��=����0���d�/����È0zE	� ��:����z�m~v�O0�ꇃ?�i��J�~����w����p��.�Z��L��,���H'lh?%�2�ԧ>��gI��;�o�����'"3�1/�ÿu?�6`��z�z��m8��y^�K���b��H�Hoyjɖ+~h����d��)�
C�*�[�u�x��}*�>�:`�#U���_rp�����-�m�;h���W�%M9�����"	o���~/0$�V>mY���p2�F%I��Hh���'�ޑV�`Pz�O]^�'������b&�6�-ut8m����}&ӕX�УS�_5N~T��?ċf��:�R�Ik2H��{j������@9�S(�t�/�dC��.�v��Q�������m�B�icA]\f_­��o�)�������F��~�*^� ������xn~���|'�$�r�����eo�L�I���ǐ��N{�{��ԓ�M�B"j��^ںMp,D�H��[��%�
=4~���!X˩I8��S�)��+��j����.�c2=:�͝q�w�O5�kҟ���`+]As}�\�9�(���q��i6"#�pf[}�}���,*+���ld����U���#�O?�j�~K��O#��z���@B��/Y�K���d�o��ph?�5�y��iA����i��Њ������4����5�&U���Y�?U�+�Ɏ:�~�Xz*A���+j��/��(��	�p���rZ�U������x��&Ll��Fs6�T���&��@�7�h\�Q�	�� ����y_�5�r�>�����e`���d������K���L���B\K��Ƥ�~5�C��)ನ@����$�?�~8��y�&�r �zz���w�0J�Щ� �����6�	���e�I�??�17	�p?B��/��p�^EE[{z>��w�9OHрav��b�p�|ք�k��0���̮R+}qV$K��}� �L�%rĈ�Y����Ń�޿���!t��"��_�[��?^���1�[���͝�֊�
I=|5�Z}�TY�X�o�r]8���o��FW�k����ԥ�j���	@Ό%ٻ������r�Ͽ ���ft9���gw�z[C֓7 ��-�G����Jk������:|P��|�Zܹ��WS�����ș��2�`�g�]�����W�5�7�|�(� r	�d�b�W_���N���l����u�e��n�"��Ow��f���e�'�y'>��	\�$�1����v�5�a�~��ױM`�\�Yظ�lR��_(��d� � w!�%��[��NW��9�2����E$Y6���Zk�n��jjD����ZN��%竇�3J^U������ٰ��'���Kw��lN���_��	��$�LQS�[��X��Dm��Nw�׾v3OLOf��J޼�}���nC��a�*طS刱���x�����Y���I�L�f��@A�x��4�C�B���.1uo�K�q�D<J�+W{~9�:(������:�}K}u�xF�`�!�9��O�Vkc:rp]/�0p��O�q�����#|�F���89�37�V5Y��,<�
ZmTZ�B� ��;�Mš��O>����e�	K��H�'�#l�oq��v�j5��YB��43�Gi�a��k���p�|��������|�hT_nݛ��]�q��}зf�Ύ��ɟ&җ����+��.��Z�[.SB�iP�.�R�62�53BI�J�Y�rw�<���r����X��~��1�9+c�M�J({d�@���
h�M���왉�z)�m��]$���ɉ3�|�d'�ٟ����s��]G�y-��Jy9��㇊_���b^�ӈɮ�N������h؅�fZ��2��ͩ�����[�]�����1�n��~��Z�u^�����={���q�p[�[�o�/�]c1�D�6�n^�,3{�!KBq�(P\�|a�BV���c5��><��0h�f�F�u��~���� |�d���ﬦ��ˍ:į��c��پ�{��P;Сs=02W�0��8�n궵�N׍�l��
>��W�y�5�`=�Nܼ�jeծT�:9���3��������x�іm�"����a��O,��fI����km|&դ�lOE�(r�镄�㥺�x9��h2��3����'M��g���y3_i�Yu����T2���t���R��#�*��	9g��\,[W)L/u���u���A��)��s���ȼ<X�0{����2��YP�"�т�.5Fr��@��.�_N�?��z��-3Wތyԡ��ܥ/�l�ݥ2Y�|�N��b	�Hhi}cz��}^����8�5�G�#��QM`�|���ea���\�
q��l�#S�#�#^�(h�����j��v��b)\Ɯϗ�M�bE��g�z{&|o�Z�d��|�'L��>�ѝ>Бw�w�rѤ�L����H�,�lQ��\�<���:��aN��m�].�xq�{�����c���(�=��2ör�>�x�������*,��ܫh��}.�/���+al!�y�X	?7d�jwyp޺��$��[ם�.j��vl_�\�9�\A�v���rQ��8���!�r���|heW'�-?f]7?`�Y�`������>eR$�
�L7����Ri���,{��a�>�l.rGP�����%�/g����؎%%e�,8�A=H�5}e�$�i�5���PNE-	Z���BB�Rel�g��Rq�*�e9��gP���f�$d�������J�6��Mf������ՀF>Tb-7����]x�X���!��r��I����=($��%p�mv�S��t�q	�\g:��IT��YcG���Zf�g�B��=�]����K�
���ҐB�r(h�c|�}Q\v����B�����Q��Lœ�r�]�����.m�z1��-����,юF�r�#Qg˥�xxy�z���([\�+6���>ƛ�S���yrN�׽��C(�5������Ꮏ�zم�^���p�v���ӆ&CA@��ؽ�t�m�PL�sRT��?�� �)�����s₝L�D��ű�+Ɣ�B?��g\O�������g���Y'�XƊ"�ߨ'����%Y�\T�SQL@cri����CCћwU+D��6x�ĭ��d,1���S�,��"�=��ܙ�W�1����}z��gէ���Q%���5���'QǘU�	2��`�{I��!:��T��Q���tO�~��)c�Pmŭ�S6�ds<<�5�c����:�z
�#Q�cy���ϣ���4���$f��5�+?X跺�Ï�gr�����?*�:�/�Q�J�b�`i�Oc�
��;�r��,�����-^�2ȑE��,�<����)r�i�>W�"�x��o��o���E��|h�>V$���$SeוhGq*�O�f?
!O,7Xm���Q|���pTp\��3�u�e��8�!��"6ጼ�v����*ά��A�.n$�*��LT�3dڃ��4Jj�������Of�<���9mc��Ԉ�����
���A*.>���0߫���"����aY�Gߧ㺉X�n�'�o��b{TO����wM]*پ�V,�m��e�S2	qٺ���®�]���#3$WܒV���B�o��g'�u�vbv�@�m�x�]���[�>"�B��"<A�o�2i�(l������t2Yl�F'�։T2�Ʊq
I%i��wZ��>�p?���u;5P���oe�m4;�Z-TfisW�==N�[i�Ze�=�]�$�)�6�$(�t�E3+��xk� ���6��e����?=@غ��|;�H�ob�`���w{N���ۊ�vfou���|5�&y8KT�Y��XN�����6�����Y�X�V18a�m˪�
Y0��?g@1e���b�T5��ʃC!�v��2�p�D|��j�~��x�vֹ�h\�~���@��/%W��Q�7��k���!.v���X�����U��nU>� V<!��S�?M&H�"�Gru2?g�����D�{�&;�,Y�n�GF�]'(���$�4�w��-��:+�\o�-��J�)w�Z0t�8X�N�+���zt��P�}N��C�����C.Ӹ�(I���;*���.���f�����"<���:\v7/M�lL�{^e1���(��E�&��S�_;�R�7
�l�
��d�jC�Vܭ���ycs�~�s	$yG��S���v��I_�1�kU``���P17�b�4o|}�c���Ѿ���6�׍m��U��`��'�g��>�,ⴼ7+橆��+�u�������H�S�p���|g=_~����Kk���kyΌ���R��x��y�:m�Tm��V�p���7�w��{��r�U���Û�����r���ƾ-c9�%�(G1[N�4*>�(��� !�{�z�t��Q����A]jY,y�C+M;s���?�dM�[ٻ�b������z�&�n�s)�n��pڼm��s���"k��\X?��w�ro<QSU�__� ݺ2>îUa�ɞj�!lu�y,Z;a�Т%���+�Y��3̺���f
ӞT�5`ܯ0(��/K��B��Y�>턞����4�I1�e�;�C7�֕�c53�uS�N�l�3��8F]{�ܭ=*�RLi'��<+�}/�Q���7���,2"�O�/��oKi'u�3����궄�6�/U�AIV'K�pY$f�&�+�hLp=�i*DD��]%�WL�צ��֧�iY~֍�kh�?�Uga�����tr#�j��	����LV[�5r�_�Zi���E������ù2Dmj�r	��p�v|!S��n7C'%Q=�/�SU�[�EݼQf�}� �8���
J��15���9��K���s2XiIv��L�RB��6��g���š��B��`�߫5/�GO_��r ʟM����[�U=m��s9�76l�@;ޕw�i�����V���F��[�n>EvPB�߇k�$�i��7�n���|�'��E���N�IO1]�ٻo��l���n=s�|�3Sԡ��~�]��V	Ңċˮ����[O7'>������O��P�?�
�B�ս���M�[����X�r���x��<�N�_�iw�(�	Hd9m�����=�a'H�1�Jq�h_o� ^yT�|`q��o�?���b�v��w��Q�).�pH�*��]���ҫR
_��J|^�ݗ>�5����17�^�����l�y���Y�1U.�P�p�?u��xGN��sy6CO�h7쓬�"4<��������)�z 
%��JO1h���2�?�!�ٝ͘�c\�"��u���Us�o�a��)�G��&Z�0�?���]٨�(��*b¡1f�G���"�X��	f�|�����"�G��B
9�z�p���%��:�Z����3g�:�
�Oʁ�x�;�h1x���� ����$��;��:M&���P�+v����W��b�L<�T�y���\�k��;��|&Fq��3M�O�:�Z��r�����ȭ�IT~DY��&`'h�))P����+}-�k�)0,���p�.����K�%����{�K�q;&�>���U��ݣ!xƶ�ې¯�&��}�A7i����M�~`�����};�W�?@cr@�r��������E��������/��R��f������;�R9��fR̭�Qe�Dj8-��~7���9L{���^��h*J'�m�G�E��CY
.�[yկ5�숨�E{*A�������4� ��Ku%c�B�	}��E�������Y���I��b��GiV
��7�J��d*�W�KO2G_��S7�˶�O�j���b�ٓN��d:j�K0Վ-���mu9R��?q}N?����=�c�9�{\�g]~S�� >��'�h��)N�y��U8����,՚+������!�3���������(q��9�t�l����mç����w���^u9
�.X-�q�ܙh�ԩ��4�&|@�o�I����{��!��)��)Z9�8��Y�/k����&A�[�ң�����qafo��.�_m��\o�[�	���G��u������b��,���ʎ�]�ǀI�߬�.q2
��D��D�t������:y��Mw���ﾛ*�S����*x+>�X��B�t�vU@���L����X�̊�
�����CFG��@�U�,����l�qp��Q�Z���s��o�Ry�X0�>W�	�� U��~�Xh9�}1%G5��|޷2���g�J�B���Ӟ��_=��i�5�6��T�\�����<���x<19>�����HF$[kQ���g�!0���?0�e	�$�H� �78zCqR��F�'n�XV���u�Q�W�q���������%�k�&{�;��ƌ©�|���#�8I�&@u�|Ά��;!
��lyo�8\�Ζ�گ�N���rВ�O��Q�y�i��Jc팪H��7Op���b�%�Y��Z�v��w�#ά&~W�n�����f_f��2�ħ�'����L��%a��s�������`=�)z4��a}��n|�[H�/ώ��"�Ŀ�����Q�$���,V'\} 
�d�J2�g��<ks�:O��Ys��H3�>��2����:Fa��#X����r�Q����^Z�Wv��t����ۦdӁ��]�u�by��`r���b\���P��f��-�[�BC��V�������U�tP�+��|Cx��6��1*�}J�H��τXV٪h1�������`d4	���r�C��=����c8�����#��l޸�@E��Mа�b�kw�4�%��.��W8�	<�T�q���Fd�9�*N�i�6�P_ߜ��5X�����4'X�g�g[�,��J��8=;ɟ�R�����KI.�
`d1�}B�ў�@3�QO;A� ��N��O$�_���p��<v	'W��2,�6�@�k#p���͢آH��4(�O��[ާ"� o8�g3���%���R�@����Θ\��af���`p[� Sp�W��G3E�Ý]���3}d\�p?	zh@�q����������.N!���f��������8�IV������z��a5�{M�	���?����ֲ�/e,�<В鶝��vBנ~�#��/NdR��@������GiA�*I	�[��cM8����غ��n��k���2�M�tۨ?_��(b �+�/��ӍHNr���ҭ������z�Z�/G�%T�xzc�b�3eL�PsF\��C�hR=F3A�)����z*��v����|h�}��� �}�C�j�fRa'P��]P��s��+,
��H���}`�et��+�3�_קn���y�gjy%?9!y�Z��=ʡB�^��Q`�m�c��l�%㏉sB���z�E(|�#IC!�izR�	�0��%�WK�Yi��W3brR��o�K,��y"S��j���ŪY�����DRJ{[�f�X8�+�TS��.�;�m�Q�p_�vSF���v���N7�,�I�2j��|9G�l`�����hϹS�b���i�F��h��=�*+PU��]J���F>C^X�2�����9S�r�U����0�	����>hG��{�`HA���VV���5���-�$Ly���L]2�Uӱ�Y(�y�cuK{HsZ�Fa���"���չMz���1MmH����� ����k+{!���tQ$$y�H #�S�O�G�]��̀�����{�|�ߝ"��[:�����I$�3�����A��n��mu
J�W���7��E���b������0�Ξ&�����<����i�r�����Y8���ۢ���i<Y��5�\����\~�T/��.�-��|�������_�q�"�p�䤥�y<��"�V���)ȕH'��⏈�E�57U�A�D���u\;ʙ쇚�ſ2��'���ԆDv&$�It�H#��cu��OL�a��˦x1E !���8�17�Jb�����Z�%S�v���M6K7��g�L'�'� �[�[�7��UP�,پ?0W^��)�P�����7�6��������J%p���G&�K� ���=������C?����Y����:�x��	/��Ga��n�"�u-�쉅\#�y���s=�h�vW'�$���x����
}����Rze��T8��3G��1�}Ѩ*�����$~R~��9�I􁚾�9z�|�:�*���>}:�=F�A� �,�1t���d�	�ʹ�"R����#��
O�v��_Ӕe;{ͫ%j�ɍ��K)ꕞy��E�@���h2�_R{��(�0iK��.�͑D��M�Q��w�^}!+����MW�^��x=T�h(�Ʃc:�q��ig�9*t[`��ML�6A�>u��8�V՗�ֿ(\���Z���4.�w��� E^��,�!Ӂ�D�ݷ�uh�Q��0���K֑�Ϥ��l��:u��y�~��Rz��wq��f�'��79�?�,���v�ҧַR�)'�Y�jC�Poy%��'�nS=�}!i2�p+8m/	�<��4$5_�qgh��<��6DHٻ���G8<����짥FVb$�X��l�S�4	��#�&���p���2��}t,����:�v ��"`I�����C�����?>���� ���}����d�n�>���+[�L�<iA�����̺�J�Z�-Q�	���`z���K���::��Y�*�cy������$����N4!�߬�m�{_����'I�n,%�$������pA���9dŃ[�*�-�6�û����Ox݈(�U�߭��
Hoͪb&ޝP��h��>��P;y���R>8�1�W6���z{�S:"�����t�%3<���0������.���$M��}�$B���>|���~������G"E�Շ��!%TmS��z���'_��<�@B0��,�)�yA`cx&	�['�[����?�f�xo�~"E�5��aV<��x��Μ�G�a�/H� �� ��*g�=XG�Kw�L<B+J[���	BxS����^ ��XOz[�Oh�Rk`r �ڬ�����M��_���H��uU�ǻ6�I+��M�onc��z��L��ڃrh��K:�q;�"���'�uw0�8̒�!��q�[��Ju>�PW�+�|����L��������l�u߂�p�
��u/Kk��x��"X9[TH�'ݘۢ	�<�:���7��0>����Q=`!�z�ͭ
�:��Y���v���<H�\j$������q��H@�9��X6~׽���] �Z7u�Okׂq�"����-������T���vˬ�6z�>�)gږ�p��[@<�v
ͱO( /I9KxN��v���ߤ'��o�թ�p5�3��H��qQT>t�!��Z&����X���-%R`�^�ګ�7?��\Dp,jy���Ʀh%�)1X���"�m@���@5��[ԤN��eD��t��y��W��Y&9
�_��a����^���6��.F�7?d-����ೌI�\^��o9K{����|
���)��_��N�r
�b�b���F�ʳO��Q�WW��B�~�:!���fl�d9�`� S�U�X��qK�^�07����@�3*! {��It1��S�)�!�!��ƿn�]}s�>����y�l�R������k��^�H���J����;8��_��(������CcX@�bM"���_ʲ&��k�I%d�?eU��ez���_��:�n�)'�XF}z��m�f�)���T���}E h�VNJ(ڻ���śX�
��2����a�{W���zW�n_��3I)�s�Kb{a���؃ �(p�T̫ޡ|��f��g�xo�,���a��=�����[��Hq�t���N��q����RC�l�0N��%���2��t�?>�(FVH�'�ɫ߂S!��I�1���:p�E�����ֽ� PZ��������帥�P����R��%ۄ�:y���@���9�E��q�~��9V�aZ��2)�'wq� ��_?���� ��Hų�unE,l�����ˤ���sp�!-1 ���W��F�����7!*�i��ߴ�%��뙜�Y񧻋�4� yF��/���������҆�@kW�På:A�vB��v��nT*�c;��Y��4�Lb�4��mܩko�S5]v�J����"?���>k�]n��0�U��0�����ؾ:������mƳ�7�>�s�����FSw[n��������vل�n=&W��V>g�Ϟo+� {����s��1�./��pkF����1��?l�<l��2-���^qTA �1U�lb��}�דes������+�k�A?Xhַ�v�/���ޘ�V>�K���Y��Ѥ �ݰb*X�=o��W�S���i$�O����Ul���x���9�Q�x>c�6�B*�7'���oDP���Mi1�J��0�L�@7Y�,�d�dxt����%˜G�0�i޷������
>"7�jD�K�����G,VX�y� 3�c���rO0�̩���q�*��#�v����6���IZI�*��r�J2�B9\�|4�z��_(��l�p|����#�MF�EȰi��P���a���FAb��ã�|���|[9�oA}́OjGq�����KN��_-�2蹗fyl	����(#��y���;�}�z�$��-�!X���9�����tMҜ�d	��¡������T��hC�����!Bo��ۊ���z?$����zCy"|ˑT6o~�����E������Z�7�g��-����۴1�dE�����zvI���EI�r���,���9�ԗ�(���W^WSr�*_�,3�-T5m��z��C�m74@ `��o�x�gI�u�x�s�W�9��;,!�2�tƢr�SYCz���`�	]v[�I�;��%�Q���D��+���cM���Bn� ����`�E�˴��"��l�5wt��|�ׇu�υ���?x���7�I��/`�b���Y�;/���|/G���J�`o{ڵ�)��W=�� /}���L�+��U��?|��G��\h%�|gse��P�:C����<0�d�����d��E��[ca�/0NO��ǌA���yAd`?L��c���L�Mn�c?��+ΐ \�0o�s0����f�z�3'�p2
'�~���'�Q^+Lv���_���֫��d8T�X.b�c�˵_k�cT��i�����E`�9Q�jR�#��u�w�4�AA��_�����;��{�8ٻ=f��'�X�y��P�nq��N��XH.�+B�U'S��ps�}�|�h~1��<M���_Ճ���`��ǩy���ܳ���N{�ln�|�剌�w����nnd�ҦUs?��z��{�k+�R� `�kޗ�	��o��;1dmB҄bt.D~'���1�H5pn���]�O���8/�lF�.=�;Z��#��<1��8�9v���9�� ڌ�,�d6��v�K�.�1���#Ϊ��s����O�BS�{����p��1�ꑄ�t�JQ��7�۞h0�!k��_e��?&d� �z�(�,�A�a6������Ю���<uFS��R2��Jn��V�?�~RG�Ni�"t��.R��j�@���ĺ.4A��7�V���گ��x�Ԫ���2�ޣ �q���Ť�|Q�ԧ?  ��'��/}��1�NS�������ixȘ��6�f	�{Pc�u�c.��/��]o��^x� ���  ��HѡM�~5^��2�{p�Wm,�n\��]�^�e*`{GD��553��^F�(<�����'�4Dl�VC&��,�vױY�5qOƧ#�:�S�@N�f$�j�x�M��0���b�	�"��$�w�N"%��Iy��gP<K�b�pe��g%�{�H
��G��͡��*��%f�q�6�MmZ$V��$n	�$�f9�(���Io���;�����-��k�.h:���'��~b��>�s�	X��c�ￜY��s�i=������;�q^�	�^2�*@�b��c�6���NҥҬ�X�G̥��v�{p�'�}2���ћ���P�����.�&<�)��+�E�oj%���>���vg��u�e��YGv�^�@��4�yN��1��W�E�9��u;����`� �L�g�s�{#a2�_���bS��KZ�з�x����^��u&��de�}�d�)CG��{ʷ?����뷍��c"; ��t5�]���ܡ+��/�>�4X�:�.'���X9��J���p��b�W����Jn�x��OeV�P����������O��y��8#����j�n��ùNeԏ('r
f'7
��._3�|s�ڝ��$&Ш��]�;�WB�)��P�{N4�|i��}���ʴQRa#�7{󻽽F����X�޵O�l��M�~:�B�Ѭ�G�}/y���x?+_�9׮�-�M&�%l�ך+�M���*c떛�~"�+��?] *�����#tg6���q��z+rl���1GiO��B��������$^ޯh]
>�Zу���\�`r)E0���z|;7��|�p�����D�xU,'z���/�����H2��`�4�v�z��`e3;t���m��#�	�u�\��:"�m�w�f��[�-_͡""��k��$�J|G�n�v9�=�}�ۊqŌG���w�>1���L�gU����RZ���	-�f��냹���Z,�wx�]��K�W�)\Ƨ�7��̖`H�����+�g ��� ����x]��:$�$ ��	�V�<��]�����}PF43��l�$�scC&�S]�d�����I���g���8m1\)8����d:xō��kgh9~
�6"��z��a��M�g,���K�0� !��S�<\	 �h�Ǵͨ��ç+8�}��������w��{�F�$-����v]��Y�mg�X��ޣ���O��8�z��9M�J2�	�O��&��.N�:�j���J"�f;��E�����eE�?��ȍ�U��˽?]��B�a:����ZW���dv��Д@;��3���X�3��q�D�?A���z	�(���ᾋ� �B���J�kypmU��KU
Ըѭ���|�9Es�
7`"eT�W�:�4n��|�=��M�٢-�u��(�h/2���}Q,-�F0x ��&���n/7r����p�$������1�^L\���nj�s�Oc�E�1��M�> "�&��P������Y4�[u�Y�/��}[���z46;�zP��/A$F����E���d($�&ch8�G���lE,
9������$͗xRJ�}�度�7��;ػǣ)u�l�}��8�L��?B�\�:��SO�-��n�g!��N�n�?����^�Kj�;�I� �5����}�����6@�|i�澉=�ðx��Po��	�7��n��M�·���p����K"i�
K�.��p�d�|&��k��aah�.\�l"c��BJ������W���'º���R�@�U;�p��M�/�%���Տ#�W
�o<�]튟c1��0�Nj�>^�� �ᇣ�A0�HR����@��hJ^��p&j��`�U�<V� !�I��S؎$5PT>�&����]�L�9��dm^U>�V0�I.7-���ÁM��K��r8�-��V�Ͱ�w����nm/8Ix�����>�z��8��o�T�f��/�p���R*�;��k�۸�Zm��/坉f��W�����%DfD����OW�D� �A��2��{]�c/����Jk���+�q��cg:d�`���`�y��k��|��I�åգ���-*M�UV�*^�Ǜ��$�s���O��9,%%�bo��%��Y�jb͗��a�=�"��^i�HF��>(��Xa�V��:�ߕ�t����B1��Y��"b:K~%+]ͣj{���Bt���� og�?lW:j�O�p�M1�K���U#E�\�z�X�:��炝�D�)Kr^9B���ԉ�@���m��j�V�=ET�� {��ҋx4:<6$���G	�g7X?Pc�T����N���#��I1]m��V���3~�9?�Z9^����w�O�/�&���^sMB��,K2#�������ޜm�q�y���iO�Ǌ��y+�P)�qqRFY�A���d���g��"ڵ��]�	�̚0��N3�4׸���&�D3E�D���sMP��+�)9׏��L����f`����r�q�;���g,~>�ʌz;��ng��q���N�Ҏ��N���h�ʸ�ƮC�>����#� �D����N�$���z�$B�@��^b�q�����6�rV�L��=����R]�=X�io��B2�&n�W��&BiI�G]��!X $��[��Qy�s�ẍ�G��oD�Ex XJ�m��W.�]z�˟雓J���`2_at��o��̳{cX��뭖���I��5��͚%��?chk~�^i�����R��a%�mq{r�<~W|Ûִ��Xv��\��=�7��^17��p/�/�<����ڸ.QUx���Bq��$�&���';�t�{�4���G��M"�Tς\b)�����mÂ�,u3*��:� y�H�ڼv�J���c9)���ވ����=C��N4	��H��_e��� ��O��Z�ݨT�dv͒�Ra_�/>��$(���)�_�?Ȁ1�':m�4���FV�}0@�9��rV��[�==�`%Aݙ�΀/�@�h��F��캵}A����Y��\~wJU��In��ʶ�Z��}���L\��"�4�ڥFیԇ��5m,���o�6x�W� &�u8��B����_O.�_|op���ąe0�i��=�F��%0�FE`mG/���+�W)TK������V~�EL�A�y�rȄ��n���]7q0X˩CS�FC�*�b�b2�����n�����vS$g+sEx�T�MD��.�������
=��/˱&��8��
(!_����l����Q�y-E���l�n��p�P��+T�Qa�2�'�=����\������"S :��ʗ��>�Hl<�4��+r�-�gU&���ΰ�s0��?��څ�_;�;m�'�v��,.��?&�6�֫�\@���Z��^���p��@����w�����_*L����Se3Ԧ#f����
������<9��!쀀���K�,!߁W�Qw+�]�Лx0�8�[*J��ݮ�>l�9�J����P{%G�a���� td���z�%���-�G��Ӟ�v0�I�����6m��=�8���h���t��w�?�:����X�K�`-ړ`N��ڝL�����q����Yt�eB��).M���h���7zC�B��^x7}R+3�14y/\z2�A\>�}r���K� ���͒�
�z��դ�QW�<V���G߃��_UNq���T�-����)���Z�A��#.�q	jǲR�2q��1ԕ�?ȧ�yO��L��Qf���t���zO���ŗ�sLgE<^vI��O���Jܓ�^�S�{��!b �@?��s�����1/�E�OC�By���C��YJ2�*t� �v+�:H%1*���E�b�o:jF{������	�|_�Ly��@"����O;l��<���T�p�+#ޛMD���)V�K+��9�Ef��6qd��@�Q�	�g�ħbM{>��H��ߧ��{�ɦ����׉i;:�39��W',L�`զ��t���$���NQ������5x���v��z��{�N7�#`�1��t�
����h��"7��@�2���p��c(DZỄ��o(�\�K�[l���G{�?��ֳ��>��pm��v�!/ �ʈ;�l@_r��%��[�23��Qy;���@t{���mq
�����j��B��Z���h�ĊWy���W8�!�O'�tq�d�bͦ��7�Sߗ�!֨Yy�ڟo��*њ��Q�/�8�q7�P�?�DHt�Xcz��:G@�$���D��k��_�z�L�9[�V2�.Th�������[��p�RBS�x�E��|�L?اC!��h����s�NLrJ�Z��̦��r@�Fb�-�=�հ0䑚��.�3������4�{q���or1;�z_�8��S�S1-K�mvw��렝�J����xu�A��`o� y����_J7G����}O� �u	n;�@V��7�ñE\���%�T�Jj�v�������[�=�>�b��3��l�DO�$Ϙ��E���v��a;��7+��^��U��urJ
�:3�J��)�۽Z=�K��)u�j�f�&�Jn�Ǌ�ܝ}o�]N/�Yƪd�.e(O��؋{vR�=�IX/T^��� Kc��ɖ��&���( m��at�_H)}ݧ`��s	���C
�M��ةA��QN[Zќ�c�2%_�ū���n��>׈J֫���8q����!���G��i&?����I7��d
\���o��S9~�u0Ӈ�U�W���{|��/W�ٮ�/�lTJz	w]u�N9NF��u� �=C��n�|����ji��ό�5V3�j�|���(��D�I����iF2�='�e�~����['�$Pou�_�v=���X`�^��-�+��}��d��I��H>�"	3�G���1�	Mo2�DYl4��>�嗂�l�z�:����<�T�WM����8�͕�&�|�����x�d�nץ�D�t����iz�1���9�"a_i�p��pɈ��z_Y�� ��p��`ӭˋ���m��#^ �H�A���QpH>��y��`6UA�	3"�ZfQ�=�LN3�n��T�����=����x����0�]7�*J}�4]eXU��I����%ݝ҈t����-%��%��]J7�p�Kw�������g�̜��Z{Ϟ1��:��\�	����"����-B�����zD�I�E���7��k�����閎���m�v�%3x�.���p׵ZZAyh>���+>�O��5�#��Om���H]�!�0����VQ+p@?E��G�L��x���#��b����dy�B!�+��fq5 TղW]oP��v-:�2S��<	x�`�|�/�&�5%����iJJ�)z_�0Ei����+NG�Ǣ[����=�+��n��Ýd#hK��+Н�Y�X��r�x�|B;@�f�G����~�YNB��iW�'qKs_Ð%�cWJ���V�Ʌ�؀'�L!������a�;��%���(0c��P
� �dKs�b�,k�0�3���@>�v���Ҏ?ʠ���Z�� ���q=2�6U��`�������0oǲ�e6��%��o4�<��X>��'>��q�V�TV���w�~�|����0�$�Zbb�I@-$ЖrU}:��Uv��U�$C4�'e���̘O`@�"#�Ļ��r��8�7�yl��q��o)�Կ���俕��ok-�(}H���q����
�5��$z�M�N��)�0�������˕s�L�h�d
������~�.@�"�\��G*�OV�V��dK��	zpR�������v����a��?��}���� �����&r�{q���f��0��=�6� �IpzM�W<{s�t\�����.���*����o%6���
x�YX�6M��XV���y��J\D��evV�ilf����@�;taҌ����;�-����m:"2�WC���	�99m�ڷ�rVϋ���eED	���t.+/�oGABZ��u��G,%����wkQL����]���:�%E?���Ee��2oc|s�,�I��c��h�l���L�$3/��p�;��R��o;_��=k�֣L6/��O���%�BM��.��=�D�F,�ć�h�#%G�.!�y�/|9��6@�Z���j�7;�O7YQ�l���~k�Ƚ��[߇8���_ݭ���P��6]�W�A�f��d��X�@�ks-f*�����hiiI��oP�D��M�?.�_^\��s	�zm�D'���<�Q_�~$�>�ϧ��N`R�NÒ�(�k�v�!�*�HQ�|��t
�Z�Y5$��«���1�s�|���~���J>��ݟ�c�qn���>,I��nֻ���S<��tY.	7�j��:Mo%8�c٭x����[�lv������c-S~�B��z_��N!�������H�/��n��]�������Q����Í&��ِgW��Cv�[��6*5�w��ݱ��|��`rj�M�5�4�%[��� W���m�~�i����pp�t�
�:�FG���T�+6X�_�	H����hW�t��$��?��V��w;oa�m+K@.�p�6�쒶��5�f	,.ϕ�߯H�����@�=S1n!��7�Hh%�V���50�˻o�~X٦��Ф�g�BO��1/"� "=i͛P�n:���آ_�`��F\TX!�?�o����^���t�)�#������&��8���c�70j�TNѮ;��:/Qь?��<m+ɫ"�n��}E��ڱs2�0�{-�kJ��d�P�߼���O�8R������nSd�{��:�C&\;4p;�W�N�����dmC$_�X,��&j1K֡M��>����s�Fvy��u��#A�_Ǿ�?��x=]-�[�㍶t�F"ܶ�z�hX�����$
5�^���#Q!H; K��������0�g�##t9��sEPjWUK>��|�0���g�ƫK��vVͤ�Q�K��� ����N���a�a��Q���m��I��7��su���[ڻϵMɔSB�Ð:w�:m��8ǐ���˖���@�|�6��v}��.�E�Sh��m���CVeU�c5y;��� ��R��t�:�ka�Aԩ���An���K��@�{�^�V�}M��{�/�Bk��9��5����E���~q"���S&~v��sy��`��U��F��:S�Nspc=����c��;�o9s_+͒��5�:��̄�(�q����٭�d�����cMol�`)��R�Q�C����j{ �y1�,P)��u.�ƥ,$�� 1S� ���5��ΰ$��7j,bQ�%���6��M���r��5U�;G<_�FѸL��Ю�6�Z���v�x�nBK�1��V����|�0�rQ}6�6&�%g|�h��$?x1QE�`e{f�k��]��R�����Ao��&����b�w��X{SW�o���92��N�Њ�'A�u��������<���
�[V�����N?��щo��7 �r��n�]�{!o���e�൙H,�|���n<Z������t=�Ē���dU �pM�;�W��s~ ��~��<Jx��(y���J_����ӣn��0X�]��RZ�Q��9���69��M�m��s�y�K�y��:���>W�tY�E�	<�x��>"T;%��a��S�����Ɏ�{��HQ]�2�x���S��v�v ������<��H�!"yZ+o`>��6fB����RLe�q�m�*m��+�.׏0YLIQbN ���sǎ�V+��M?>�8�C��=?���ү-�~'pA�$'Qی��쩂GoJtF�걞t-3������;4[M���z�*.�����Lr�[��3�x᠉{�Y5��G�ׁb��λ�_�Nῒ�-������|�6�5x4�	jG�(���r
����@Edņ*Xy�MONsw�\��`���nX=F�I[e��E$��:~f�Z��]I��4zϛ��#ō򪮁���O�8��3V�̆v�����=�pZ]����WMq"��r9c*�v��j�����N�k��/v'$7�ʫj|��2R�bm�����V�>���A~��<=�����)�����cv�/�B4��lT��!#V0+v�œcGM&��
���A�)!ǐHzs9���>/7!T�4w)��H�m�N�Y;����Q�����Z�ё����O��� ����c�hHl�f)d�XM9/8��ӵ)�{���V��Y�����EnZ�����i&J�1g�UR�7+mN�.�Td)!>p�d�qĸ���������x#��Q��ߛ�����%CНK���_s� د��ە��t�Ba��\� �*2s�R	ސ��ɧ��ܩ��LRon�S�C"�e�x�i�ݘ�Z
��n�����4U�|��� mH���I���1dc�)�x��/e�r�wj��Z+ͼ��VX�k.KU�{�Ϝ�=��/���/�;��Q?z�h�"�0~Wx��K�!~0˄�z���aU&^}�5�Z&U��j�C*�~R�z8�i%a���91��Ƽ�6"����r<@#���Y��Zlv�_������?(�;>yy,�Iw���yȬ���$�=Ǡ�j���1�UVT�XǤ;��"pҼ]VE��)	+����yڙ��g:2JO���r �n��dj�;þ���s�-N��`W:�f�աPȊ�u�D�:�qX$q_�#�~��\��+����#���u+]�2?��	�(��}߹�h�;��\����p��0�$8�&"�|��^PyӰȾC�R�ZA�WE�(�C�(V�E���h|H� K��r�ä/l	z�%��������[Z������T,�ܺI�1&���k@Z��{�a��Tcq#}���(�WeJP�ň�D-H���/�	6K!�6��_4�5�E�5�>��� [v&����[X��"��� ��º0���e��p���d�uթ;��yK*�y硆F�EY�ն+�,�� �g�|+��^yD���>�ǀ'PYP\]�m�2�*8D�r��n��ߜ�����w���7�W�`�-_a� @*ɱ� �:�����n�5}�)ZZmq��38��SԲ�v˟�p��Jb
k��:ߚ}�mE"�N�̔Z���2Z༙���(�V$�)<��c�\�v٦*�u�ȏ�K�|��"��r7�p@Ax�镇U9��6�ճ5���<yIbج�3�*���^��-c����� ��-lʥ�=��Uhz��1��S;�5BW�T��]���``p�� ���\Г���2V4���yNV۟�UL���$�U�� aB���:�e���az؞�$��dϸ<W������͡hXw�.1�yN�aiV��]'�"O�jZ�ɸ'����F�!f�s{�J�k$�PvY#[���h���@�9B��$M��;+=�$.ǃRѫO���/�����;��Fӯ⑱香|��~���&a� 
�����'A�w��A��y��i\�|��cæF��$�x *\N�|�j�WL���@�n	ш�㢓A�����{>�6W�ߗ�]
:#@��7�#ix��F����lS3���}C�P��Qa��!�v��l�\9B*�*!�jV|N�єF
3��ʬ��G�&a�k���":�'�ǁ�B���Oz�
-r�&�bi�7���������T)�O���������s���V�7OQ�Ue��O�����9��"R@������'�����	\V�O�VZɮG�D�O{پ�����IF�J�-M�S�a��������*�!���(~+�1�c�ݞ�7k���6w�!V�7cT��Sh:|4;�ɨ�1G��b5�=��#Z�BE��ϕ§�r�|�p�h|��xU��p��z��z&��*�r*������93����]k�C9�C\���v�跧r�:�� �����݇w�P�����n���ÃW�_��/�c���?!��[�=��us��<�~Sd�{c#��1h��D�=����?���N�����v�-��c�J�{i��@P-�l�U�a��}�! ]������w{M���ir�5fG���3>^5��ļw�aNH�0J�����X�%�&�N_�In�, ����2��\�v4v�e��bg��I�Cq�������@j��!��d�/���������,�R��
Oꅾ����P}�B���� m�����-�t�"z6!����Ht9<�����U��N߇$*��؟���:�^�Z��!����YI��w�v��(6��sUF>����߹�e>�I��UlF0x9�cL�w��;(��\)�U ?Q P�z�/��kE�e=�C��e�R��t���ڛ7x�s���"���!�>N�zm��:�{�VG��/�����Y��5nW89g~�-���2������vz*ռ��BC��(;�O�:��U��W�!Q$D�yEv?�k(��_1��'3��"���F�	��ѹu{���;w���u�W4Y-L����6��c��-�< �[��*t�b�g���6k���Yu��t�f�6���䌼����;l�O������f-�L�'�K;�%�Кm��]�M~C���ӌ��]��g�0>��v�[����j����h�z�摦9^z�n� A�·��1���9v�Ym�_�9��J� ��x�2�#A��G�}����u������fl/��.���4���lD�
Qahv�������X��!
�t�}�1.-��IZ�� �Hő
[G�⺙�I�yT!O�_sQ��qI+D�e�!�>���gtțQ�\G��t;Z4�9��'t��DF��K���N��/X;�B�_Eo?���Y��w^��&����)��J�;�F{א��y��-���_�H�n6xe�;s]��6 ��B�s;���֫M�E�G>u�.R���w���7���?w9�%ī7T��IhЕٞ�P��s��x:3ԟ��^3=~��`� �H�v��nN�Y��7����Җ���(����&S"^��[�Å���U�σՎ�,R)w���CT|b�ߌ}x��7l,�F�7�'gɮ��()����峆��ʀ��� 0�Lv�ㆅ�Ў�!�bk/?��0X�_#x��D{�L\!���:��Y�T�z����a�ކn�*�u���5d�!Vm����r�+�5�5����FW�Q�*�jo$"G�$��+V��S�ק�o�VJ}ao���6�-'3?'ҩ4Ɖ�Kݑ���H(��ؠ�ܾ�{�v���i 3�'�۷5ew��kn�@���	�&����z�
�c�r��'�p��`�HxY���6����̫I�Sch��-����X�3�����3��A�m�& �u�cFͺHty�o��No5���j�BU|���v擥p���5 !KҠS�t�~C�$q�ũ��'���������m�=��U��? U��r_7�%q��[�7j?�V�Z�0�`&�9�a�w���'��T5_fq}�a��1&o�ڤ��.<�g� .��ߘ��>;Щcύ�z����e)��Z�s��8ě?���� ^��EFK�m/��4�]�zA6<�Y_9G�]�2$Py��>�HsR8��d
"~��]������*��������7���E�}�x�mjt�Q�e��
��lغ�+��˨ ��v��g؇��u"�Zir���G�mqOr?�Tz�EXe�#"t�^.5�.�~�	0�A���9��v|>�<��?�ɾ����M�o/��?���d��h���Lg/?��Q�q�CE��� h=�qYy%�ڲ\n*���[B�C���IH 2i�6���ɮ*���>$���ݿK"�DN'����f�5��u��Pn�Zo�ᚱ�tK �lWM�S�<:���\p������!�L�|�?�G+�m,;�o��������l�Z���䁆��o}nOu����-����ȞZtb-R���/7�O�d4�K��	�;6�V�f����ZE��D�ˏ�j?�8�x~Ȣ�#��۶�T)|>L�]B�!ⲧ����l���_X���(�OlW�ֲ�$�S�4��ٷ�%U�$$(*���VZLYc5��貯^�ؑ��
_P����:9�w�Y�v ��rvOs���/e�+MH��Fa��,�ڿ�.fp)�
^�h��#�F�����Pk�"���{�����A�,U��e�kd���� ��J��M��}�vw'��Xw�\��%#B��m��>	��ٺ��7��ɱ��*Uu��{���w�I�m����3��_�QM�����r^�$�6��ɿ�mt�̀���@.��D�	�|�uK���sR0�#1 �v+��ro���S�}(�Ӭ}>V6���l���{�IO��Y�Ec��5�;7�b��[�J_N���h�Q�~�!���]�k�A~��$��*bz�)�yas,��>���"��
�u��!���d��ӡh3.�I�2$n|N뷝�l�X*B�>䗕��A��|�� ����v�ӊp2��׋f�!�hO�mh�{�vk���&o	=LwN��yㅞ����*����j,�4�w�M�H�)�(.B�����l��-��"6�R9k��i�nI�}�;��U~q�X�4΅�%
�C3�%Ch�1���Aw�m��D{����,��Pc6�E��yn~��
 iDm�A��r��HEݔ���>�Jc��Pަ�Tt���,A7�,�Ph���t�Ƅ'�	�<>�����	�D�J�ȏ�8�{h�1�|�g@�l�R��3r+��P����B���WS�X�=<߫��.3��G�V��(y
�;�/�݄EZKݼ��7��
��3�SNƖ���T��8ݗ�3X��q:'��̥>�ROgj��9�aV����
[�%��(i����DףE�Y���-b�W�C+���{�G\��M�C@j���?ȧ���_���Ҍ�-o}�D&l���Rm��TÖ�=,�nkO�O(m�V���{"�Os�F�������4cn��CZ������K^޽������Zʺ���^Q;B�R���P�Գp��&��Y��@؄H������?m��� x7��\#j�<�^�b�}�H<���Ｋ�?��s?�+��g��K�Oӹ��2�|!V6C�Rh��JtW��YG`I�\��\h��'Q�~��yT�O�c���W�p��p��r�j���XN��n
 ��?#��C�ɟ�8�ũ��V���ř�CR;b�/�۱c��Gر<��f��u�=���S��~Æ8y�~M�h�H�;�a%�:���3J����-������GІ�/�0��T�T��Ped�2=�4#�rX��;���v����� q_�VRh���3�F'����}E��b����T̙7O��Mb���0�u�))	���?}\_]j'"t�sƘ!|���e��wX��k�]NWw'�''y�~�C�y\4�,J�L��P$��Y�Z�0�C���G��,����m$�����z������%���-�<�Wk�RmJ^���t�}���X�D��K[�,򄝇�?��_�$+�f5"�?|͕�w��bIPc��e�C�o�bM����:��_qg\�����;�����ꗉ6:��i�"�[-_F+N�n��������}�;���5�X�=f[% ��G���6��śk�-P���#a��Y-�����a8&��Y)P��H�/��C�q�K���a�V0S>�ԥ)�L�2�>��M�a\� ���{����l �yV��z�����0q���-�����9a�p�V#�?B�Ԡ��Y+�_y������w�M�	\��&���45�,3�=�#A�wP�"�~���ɺ���:����
p���F�5�s(2�H����{��%�� ݤ8+N�("�Q�t����"R����<`1��P�J�G�a�?��U��X&\�s�w����������؈�i�o����/ 4�R��@�-q�m�榐�N�_��]ޠ�Ǐ�:��z[�?�{�5�����mF��|�m�66ޱH
ʮ֏d����ʵ�X�v�JZ)'�����{zi?[̙Ԃ�.�t���z�4B/���B'��d���]�$�(Tb��w)R�j��"�F�;M{ۣ�xZ]J=�6��F@�x���gGĵ���R�Ngca?|R�2���w1߄ _8��\����Z0Z�^�CeC�ݏA$���R�L�"	�@>�V֯�:�RN&JX��h!〸��ǳ���c����x��ڙ��(����r�Gt\�V��$�w��2v�w���YƤνǼ���)�7���s��e�-�(�����ݎj� �Y��zd�wr�X���v3�,"�r����Q�X��.���%A���L6��G�nh��C��?��納�����*���j�������ԕ����̯8�)�T,qM�A�c),�*�,���^ �)�ܩ{�MZ�l���d~���Ȏ�ć�?�! ���g���-�-�����U���2�OD�D2�M������o���݄�/ߤ*��C�ho}:��_�p�փ%$������P%J�|�	\)Б.��\���H:����~7�����j$��6Ar���c�$�$z���Q�<_Y럜�� ?�)M|�ۖ�O�����m֪Fßi7����A%[���'e��'�-Y4T�q�;n���8N	ߤ��j)V FJ��wU�!K}�G�n�lf�R����aW�������/�!A���c��k�l�onD��Y����;O��m��+����nl��5#s��c�q�?��YM��'�l�s	�z9V�)i���!b֏�J�Ɯ��ZSxc��;�F�WK>AH�ג�3�Y��b�kM�K����X�u�X������<�1� �4�dQU���H7�է�\	j!)4��z̟��_�)`0'��fU@����] >����8��������}�Vｈ�"�?�W,\�$�&m�kFm��b.ޛr6�����*8��(A�wX�t1�8��#���x}��q,�������pr�)����0��o=��C¢5��W�dط���Fި}������!�b�]�K7�ە���Θ�
� �7|	0��"7��=��E�*~B�)����N� �p��v��*V=��-�ٿ:oz����}| T�ᯭ��h�i��_�!�+��jO�^�����m���? R����q��@����;���Rک���^�EGZ���#{3�qڴ��_�L�.�<"��s�
ߍN�+�\Ȣ��X�@�rܻ�*�\��?0�4,�&�Ї��k�l��Ñ��;_�^3�-��V��`Vt��}��sv�;"��*��򫃹�I�H?���.^y(�p-�'b�E`����;�
Ԅ4[0��Ms%Ѳ@��������-�Ј�b�J���x�!���Z��.�E�R>����Gy2�����,�7!��B�K�E�4N�<�}� w1��Tm�E�j��)�5�:�se�7ϫ��4D�$\�Ys ��X��K��4I���pEñmK��ǚ�$�Zs�=)�}�ɦ��r���u�#ߘ3nJ^>
ч���J#��P��n�C�w�Wۡ��nz%g�~�l���S�6@<0d�b�A[�)�ETW�Tn+��+����y��C+���]<�rgӪ��ł�liB�. �Z3��yܔ��W(���[�!�u�t������F�V�.E����gZ ���Ƿ~P�f+Sέ&���O���R���}M��Tܾ��r��W��^e%���21
�u4(�2�t�^�2Ju)�Y��-]��Xu��]R��+�D)Ua�F�7�f�����-N5�)}-�B[���:l�ٟ*������zD|�� ���Ӱ(�W���T�z���β쿊d�V'ʋ �1��3Q�u%J��=YO����<�(� ��hJl	��-��X�����	yX)֪փ2զ#:ѻH 2�튔����Tg����c{��N��ʛ�1{Z�J*U��f�Q�%� >���ڝqtA��c>�9V����E�M����K������l��b��-�|�D<m/���Q��:���f�dز
�[%�us�hX�Z�h�i�X���"�����tx�i,��������d�ҭR�2����~��p`�)�i`)/�x��6F��7O�o���+���tkn[��1��q��5@�������y��Į�CL�gj�Y�7���q\�z�*��&���sD\��\�s�+I)2R�l�:����f�z=\w�Ki�yk���¹���HX%�ԃx�m�M�(Ch�^h�/zU�Bd��T-U��bO���Na��߹��y�1{;������ߡ��9A�ûi�S�3T:��Ʉ5�L�y��7
�:��)�pG�I(	1���M<߹���4L��?J�r"����ܕ}�:u�sM��t&�S�����>�o���2���1 !N:^����cl�_;�(�����!�oT��b��n�镢�^y )���A���/�q(��I��9�?ƩDz�"�n�<IFB;>����ؙ��K���t�g��_����vxق�a���G)%o�\G���ɧ�i���$v}�j-�Y�ǭsQ�����wԒ��B����bh�����
^ˎT���&�-�}��3�	�q/�c :$G�ָC3��bS����37�H�#������J ���g��
\	D�+G�Q1�:Q���;��� ��"�?��|x�S�&{Tf� �2R\�G&��cq�q�⡏.��~	��\����2�7v�
�Hj��,�ŗ�x��2YO�
t�TP��	^ZҢB]�f�o*)S%K`�3��m�d*[��!��|#,}?`� <��>�}��c���U�!-#�jc�_dhS{@)�T�f�q�!r��]�R�p4NA��3 �BБ�'Bt|vū�=���x��jGS�����e[=u+?���~�wq���>�b~8|��7Y#�gpr�4Jƫ ^�6�%Y�><��6�j��9�Jt����/����{��Ul�"&%Q�5b'
�����V��Ia�"��'<w�hFa������OxC�_��/�La��Pq��\���ט�>Ƹ؝�s�=�ktܖF����IS����^y��o�I�Kn�Ӑ���Y��:V��?��*�J��Ѹ#(���/5�m�4�����������+�}w_;XY=]-�����XB�=a�˒3�y�D�߄�4�&|�msY�����rA~h3�l>Xh�x���3ɷ�
U:��w�|h�,�c���q�0�d�S=�>�6-�"��zF����J�g��ȳF�Y{�0�U�X����[�,��C��yc�jQ��c>x���Hmq�$�B��E#�)���	��H��c�T_�S��̡�u�.��$:*���r;��p6��;�.�h|�A��4�[z �ςk�c��e�:F���}q�)+�r��
�b�9H��;E��`s��=�����yz<����������{����T,'�w�ϖ�8=E�k�e�[A��r�� t�K�
�3,e��C�9�4�;xC�K���OI?����'9�,��ґ���u��V���
n�{�n~a5�m��>E���ouҡ_1��(�x�@;�l?��h��Ƕzg,՛���!����3��K�t�b�-�4S�ƛl`BI�B�>"A��;�`��5b
��9�Dْ퀓g� ������nf�0��!�6k�A"��ړ�6�P0������BU��T37��{D�#AM�
ÎV�L��(��=x�;e���4s�#h��,8���B���*#Q��xv����&m�p���g5[eP0�"��r��ΈS-��!�]<S��V�^��ح,k,
��P�:��<����)!���I�f��f�g�k.ud1���̵ ��D]{�����Mm�`�&�9��XD��#a7��zR���'�������/V�������GP��6+:�k(
^�L���-]9�qժu�l��cN��)$��CE5��7i���xh#�[(������Y{O����'�jߧ:���%	/��ޖ��w�#��Ut>�sM-Z�|8tS�Jz�%��~���O{4���g��GuS��J��S��K]��Qp?�x�����~��}*�n��d�?��Փ1��3 5���JЪd�����)A�P��W� '�V����s�h	�#��:>�lgG�JQ�r �s�D���N�:� �2w۷��-����+P�����2��,����[�3}w%�C�i��8#\���fU�A���˂U6o9٬6��hP�$)QG�v�>�u
SU@PEEy�����UWf�}��gue�'�IHZ�c)���!�Ua��eE�<~ᛧ����P�Z@��
/�6B3�s^��;�0�Z�R�řN
1:��҄<k���@{��\1d*��wh0�45�R���I߀�Ӄğ���oX������@��S#y����o���}nY��q������ɮ��p_�ܭ��U�,�BZ�Ì����qC��/S;g�\�y]
�B�)^L�U�\�mk�%KwF��Ȗɞ�MM�ZM	]��YWz�������3��JZ�^�м��_���J'VG�dWbuA@�$t[$rh7Xs�5���.�$I;Y}�x��
0Ұ¦|K�?��Z�D����&��V�6���׾T����b޶�:����A�0Gۥ~�.�h����RC�JzҴ�������<Lr�@♷�f(S(�I+~��rW�_��MG^�.�=O#)W��}!�p�0�I��Fh�C��wDt�I���>�%h��O�؈y6�W�--�d:܋�����W���W�j�|b��\�j(��x��vG��7%��qz�,���yn !T��D�Uo�]#��
�~9bEh|�f>o��5ve��7����U��9��dQ�E{�r��-�BE>������F-M�Z��?�9�>D�p5i�"�B��O:,�#��;���H���
�K��!��&3���!�\9wJ������XO���Yx�=��h�-/#����[���Bg���4V��H��R�e�H�$eB��O4��9�=SG�{
�uv7uū����9����hJFA'|�x0F�kb�d\�ߪU���a�%���ֺ#@wA���K��!
�YE����X��>�X���S^����������#^���u�[�tL��>-7z]�u|��wN�T���rx]�M�x�{�-:��mvx�v�d��Μ֗��{��r`�E��s�#�+Ǝi����w��rӵe�����g؎��VY4S?�x�~�	�F"P�n9o'x}P^�8Q��q�{Az�2�oJ�rB}T���֞Ǟ�絞
��c� �X��^e������2�L`m���	<¶�����uxs�ѱ���z�E��:���~��I���Ih�[PO0��҅��:W����A]�'^˘��7DT��.���y>����տ���%_q��d��G��*�/�T��?Ż-�=����‌�!!%�;Z���ώ�+���s��F���*�O���q[i+$�;�X�yT!�L��T4uy�s��d��1����-C>z��43�7rG�X��&�!���3�"S*�;
�䤂N�jg�d�ί5%�R��+t�-f��3)���@���݇H����D[�5��!b�]�3�I��sN^���c�tj�#S{&e���o�yc��aI�b�]q�j  �$S��W)M�Z�T�n<�C����[H�0׆40U44�S*8b�� 2>���l<��f�������d�Bo_������FA����z��w#*��1{襡�,5~7zk��KJ�
�3����n޽%��Z�="A\���[��&�Å��0��97�ZT��[�9�z_������z��߮�������v�E(�Nf�\��4���ew��֑��;ɞ�oe5?��G	�3<�O�&���9��x�Ҝ=<0���>X�1�{l�	�4'����K|���!���h��ZH�4����
�a/�$���ȧ-�xő�Z�1SOwq��8�2���+���e�H"
��3�-|�T�8����'�SyUg���4h�fL0��h��	���Q�����KQ�x	�^Z0����"lw��ݝlP2a�WhM�K^�@E@���
6�w���K� y	���!)���C�0?s��qn���#:w�v�p�ߗt$3�x����B9-}��=�S�������)�t9Â���Q͐��Y�2�k�1`��>�cQ䞣Z��C$��o|k�6����s�4�M�i�Ư(�c�A9,m�~����܏v�W�煪�
�m�y�@zA�U�FS��)��������]�#� !�����`�%H��y�bx��t#��,�����~��q��.r8/Q�8N��
�/ z2��p�l����YT!&�q
�&f���~�Ԙ����^���b����V�0��1U8�@��i��!7�@GF5��m6ծ�~6���/F�B�"�t�W��_]��s^ci�mOZ���
�>mn�齘=���qߐ����c1���,�'��,K�;�ںG�D�o���>K�0]h�nW��m��imF�!��L������3�d��|d��>�<��
�%��7�?�-^�SXB�D��'-i��7p����䏞�GxX�6�[�L����.�T�
Q�|�2oW�6H�7�����>��Ic�fl<�+y!?�-z�la"�_��c�ߓ�h]�TR:��	�6�&|�6i�qr����lNr��¥�i/>Ƨ??=hO�u;��-���L�n0��[5��m~q�(������t �e�K�~w8]��`�H9	��C�O�I�pR��,_���(Z��<$�{+h#�����$Y����*kh���P�?w�M_�[E�h�$5�q�~��B���㴘r�З j?�
�kf���袋}1���ǳ����T�ri5���C���C<c�KO_�ZMH(�k���o�S�e��ũ��vH�qž�����G��U�Z/��Uݚ�R6���NbШ�6�����)i73�T�A׊-��6h���3�Ti�=iL:��&��4ݷ�*���Wd�e���^"�A�"H�����m	9�WC3m�l���Ɲ23e���/�;;���{��1�`1+���0m^�҆8��}�g�famu�v�%�>�]��{y�lc�G���p���/�ɥ�|̺����#f��1�/Oqǧ*�h�iuR;�.�h]O�K��3���X=�G�w�{{mQ�"yW��rw&��Q�`N��x��`���r��<\�P��@�����|$�����FQ�ϊ�~�B�����K�זˋ9��������/<ܭ�F����}F�o�Z�)�6HS��ױ؆͓���MG#])�e0��+��η�ؼ�O�%���_�[e{�w\}`B�k<#��d�D�.S�B��7�͎nj�v�F�f��-��b�5�������ʑ�Ouk��T2^M�i��MTQ&`'�z�A@9�7���%�1�e�'ﶝ�3��ì*���p�����nw�r};S�~�Т���$��z��*�d�~��wk�n���رv�}2��DA@���\�w��ѯ�A���5t*�m���Tj�$�����ڜ������$G��,/f�Hx�2{������@�Iz��)�G�g��ߠH�ðVn��M������o����t�r��D3�ܩl�7���q����m��U9��3�^w���UU~f����f��2fH!�l���n�yw�C[�dy�7�x���<C[�a� 4� ��}z���Z��ߴ��!b�6�� ��T�#2�Lջ� S�~��մ��O�ê�K���1��v��7_2��Y�ͽ��~Q?�:�K�iQ�/���n�/R��:-Q�oO83��W<Y~��Ae��
�y��@� 4��X�v!����I7MB�������mP�u���D)�&��__�ͭ+��~O^Xa�t`Q)�.��J%����Mv�{)�q�=ay��c�*���n��P�[��Ŋ���Nq+�ݡ@q/��������K�"�|��~����M���{��3�6RV��^t@�.����ۖ�T��cU�` �Sk��-�+<���p�1.�q)H(͍��&�D4���=!���J���4�*B0�!l�,�G)؏��jp҇���WT��X��b�E��qq^4�i���^dh��� �������\Q$(3�I�ͱ�$q��@�cI�|&��YYjі����X3��o�fO�kk�X�����2���j��X{R-�@�DCי�/�>6��>dj�xsZo���
-&K�Z�O���q�.j�/Dy�S���3*O�F$w�Vf����[!�������r��Q��I�X�L�^I���ӫOf�U��:�?$�l�+�=���D�$���&ɹL�7�O���11��<���Oɽ;І%T�Ȏ�Zx��g ]�]Ώ��ezB/�(�:��K,���'d��ȭ�2��v�CrIn�	���0����v#��e��ʏ�,Є�M�
?��֐�ow�U�-��H.VA�=O吏L3O�'�1���v���l�f��/��,�@�S )s���iʛ�㭋��"��"�]*&v�F�����0�Q����1�51cm�u;���ֿ�;��=D�^��~��ݗv9�}�1�K�2/�
�u��dE7v!�����Ϫ�
�-@u�qz����~�Hʨ�ke]��BD~RiN��H�"���p�x��y��(�&�5+��V��ʙ(������I����p��O�C�&1⫔�J0�J���vS'g��w�a����_������3�;o�[�e4xHiQ�~|�|M����Pm����Ku=[����"^2I��˃Ŏ�2�H{΢�`��y�F��ʩ9٬�(TB��um��y��U���=kL6��E��%���>����P��8���w�x�+�}* ,_��ߤ��.�{3��oX&T|䁨(����ɟR�f���A�`�g2���]��GJ�=�^2�����n�n~!#���9�ڭ�i�H\�%�����[?֢>Q��K?ՏRd�-��N��6 4N�h���= ��Q����|��'����������ﱔ�o�C����C��xb�fK�X�`7��BŝRl�P�k�o��z��?�|���GM��S����>���Eŧ'ñ�_�fT`&�E���"��%�5�گ���D�Gx��NU�YI�?����I��+k��Us]���J�ŏ�gh+)G~4�Ʊ����v14��\ƶCA�]+���
�����d>��J����g�_�Y�PЙ&>s�N���8s�΄�0Ǳ��^h�}}�N���aJ�%���h��҃�g�����r�W��%EBP3�k��/X���kS�4�Ty��ٜ�cS��z��͆�s�	���N��.��!H�#���|Z�$J_!I
9v6J�:*��Kø�j�#��Z��_�̏'Ǯ�aP)��M�O��u���G�#��kc��ä*�8�ɑX����Y.�2���ێQ��G�#I���Ȉ���k��&�*gx_�ć�)j~>N�yRqBWxֵ�,�-�߅����k�'y>��)����
!8s�O�k�QB�M����]����Ӗ��F/|`��"x~�2�T��23�]:J����/^�<3�|�ʉ�`-��D������N���8�"��'	DD�0K�gq�:˦��o9}�Y�k�\4��gqf���P�8kaC�RW��ca�lJ܃CM;0���s�P�b��"A>0���=)��&��t]w@H�rҸ	vtmMވ���qa�ͤ
�vWѡ�������(��%����镤�A�����q�*�(����U7u�\����̰�0D���bb?a�j6G��1d�کY@u;����u_]���'hp��2nEn�7q��-�TZ-�x�o��M!��15�)���p}�ݏ$i�VU�@��z��6���UDz�2'j ��z�/��4D�OH��:%�`�~�8�@Y}
Z �����D�{�Q�c8���w9�

���������$��R�h!|Pn1�X��{|JEa�~����O�,�½�z��mZ�ظʹJ������h���\k�^�^r{��'��"RJ桧�����@��g+G)�P�s����HFЩ����THF]&k&T!����n�4��sD;�*9I��_*���i��BU���_Z�ťц�{�y�pξwLu�t�����Y�
��T����|�z�}���d�~�=��u�u�.z�.a��?��E���L��t�Mx�h��v=�C�iZ#�Tfr������n�!��	qg\)[�Ԏ�{b���	0�߃yJ��{y�*�[�?#�i�W�9pN�dݥC�)��j���)���^s�p�}����e9U>׭�ԝ��yk=쿖�m��P�8���_ӓ�������fq�i���z�u����:���&�c���+@"�=�[�������0_Q�i� ��M�^L2>�%�?)�í��jT`>_���W���U�",cR��8֮?����τ���9j��5�S������Z��P����<"�H<ΙZF�<�<�3��G=��esn(h���e�*� o%]��_�$FG�6�b����{�=뽸0 �V�͑$���=����G�,ֆ�j�i�Bq���!�Wj���?Cѐ��sQD��V����&ߞ?��T�r[�g�oX�I���A���[|K`Nլ���N
c5-r}Z���%0C���pK�@쟻�	��ze~�sGhy3��Ԩ�!Eê�S��i��g�Q����Ќ�7������|�C�� ��Ɖ�(>��E�D���89�-�s�5����!2|0�}���.�>�$���;A�Շx-2���F�+E���������^�v���ۺ0o[���=�,)�ǎg�ہA��[�����8���,�pd��	.�!�|�_��$��Od��))|���a�ȝؓqk��A*� ���8{��rs���(��Y�X����Zt�h�ˍ��8�{Yp۱v-�t��
- �tn1T�����01˸�㢀�!�w�O��%�u������7b
�|�~�o�� ��B��0
���]�{�￐��f�����C��L6�9I]i~G=�),�8�3���Z�I2y���a�P����$��� �����Qw�~�o�c�Mk{<��:c�it���G��h�[�k�����[�*�߯`.(�v�~��:������"x���(��גw����g�]ؼG�K����8�5A9�+��֏m��j]X�1�7ZT��P,߼��jV�}��ylK�{o��>�{%/�u3ǽe�D|z�����ll�������Di�h��mY�4�4��Z�3����e���rǻ���O_��}��~����bM�`��p6�@�n��M{Ar|���{�� �R����D`���V^�7"ʈ��C������=�o��x�AX�n�2�L��܋+a50���,5����[.�D���L?�c*�����6�����k����=�07�<��9W�K��z�ͪ����M	,�׳w�o���d��s��2�� q^mϣu6�ߜ8��3�xϬ��w���f���t0*^|guٲ&��D�ѳ/���0��ކG�܋��&uɞ�$��e�UT����{��PO^�}V������W[ޅaO*%���7�	� zw܌d�yB�z�B�#9��EaI.�%x����C"|��~�������j�Y1o)@��m>3��8P��T"!�6R't(n���S�l"|�<Tۻ�#~���:����>��"ѭ5�F+IS�Ds����B�HF5#�_u��܈[�oT)F�q��m,�Ь�p0���H�/~�HY��#��#�^j��n��-� �	��l�8R`���=qN�q���֚��1�ߏ�k�@��U6�����̷R6}���E�A�R3�z���Wx�I�A����qɩ~�rE��{����
��֦ga�7(=�B.S��+<�S{<e�39`v�'�c���Q�u�������`g���|V�M����F�Ӛ�R�@��x�B��6[�!��}�����I�i��l%�Y�ܗ��Q.7��cX��[&|8G�1�T�
P-@�NƇ����_����h���9g�a���4D?`�d�Yo�L�h.p�pˮ~�\��Y�߂��k�o[�V��w���V��\)ی�Qe�窚����\�Y�����lB��&q�VF�%�1��ʒ"V[v�n Ǩ���J&��B���e�<�[�Q�Fьb�u������;"g#ec���S6վ�'LCO�_�CT�7��>�ZN��\ߎ�xىTB���]�Mi�����%]��RqcJ�}Qv��!u�����G��!����2j��rm}7!wӍ�x����F�!]ϝ��gY�˹0�H-G��]}��#l�=��5��K~K�y�y��Խ�'WLZE�G�YT"��� �/If�M��pe/�Rk�u�Ѵd��n��z������$O�h�>�k��*��-��UV�C�
h7�������y������C��U��߾�Co:C?�g<�n,}��H*�WB=u�9�,�˴�����ڛ�瀨�#+u����q�CC�@��-����i89�q��$k����n�/��Rf��o���j\p�F���j !��˝�:��Gb�u�x�y�EV����P:���Zz�"��e�	�0=�P�<�Z9.<5�E�L�a��<�����r����u �-�ml���T0a	���'?h��V>�6`��p�i�� Re^4�X�g�{�X�����p�w���p���@����J��K�����=.����* |,h.�r-!�σ�<��P�P� �EnD��J����nュ�¼NeW����}x=(��^g�&įY�9]����:��8���?�rك�4������a~*�t�*a�!V�?�n��D�u��.���>��8�*p���z4�bߴ�1\s36���P�O>��Sү]�"o<�Q]��W�"O�B��U�Yo��$�(��4ɪ�쒤¯�ɣ�nOӂK_b��l#+�<9��,oI�.%7�r�ɛ�n��O��(|�j�L��0�x������!A@�[�b������!�p�����)�0����z~�=0�Q�.�m�J�Y!u�);�)��%<� ��CM�_�w��\�N�{�OG����cfa�Lvc�6{ǂ!���m�O��M�J�+T���o��>=ބ�Ҹ^6~�>�5eK�û�3 B�g@סt�S��#�'�� j�B-0m�g�Ut�c�D�Dr)�w�α�o��;2\��a�y"c`��c]l	F���d{B^<��\&E�ೱ�yC1�<'Kˠ|���J����e��$=T�ȅ�zS#0�I�D����~�O濇Vj+>_G/ӑ����8��'���=�����˪S�Ŵ%IDS��p\�uGfP����2����Մp�;��U�T���>�[~~�e�7w�~��:ҵ?s\rU(:��2O,�l�H%L�����iM� �t�j�ؔ��9�RPB��+�V��lE����W(�c�)�x��]����m����d�4��0��Bm����Ѻ�"�g?��$V֠�>��BѶ���}���3����xx:� ����3κi�Q.����u�B�U���[~I�t�zb����E����S���jH���_bޘ��_x�(�W�j�H�@l�cb����չ8>�s���X�/�BO�n�y��Z�����!/据�tL�ez��������x3�1_���4�	*_*�c��n/w	{�-!�ǻv� @�4#(��ô"�?[ª�ByU��U��+��h���.� V�p0r4/M�|+�p�	+��[�J���8ξ�L��q� 2�9�Y���Co�4O��=����ƿ@I�I�ql%�!�l��9��Y��k[��Hx��i�J�����&!�Z��]�u!d��NT���[�ھ�|��3:T��%v���N׌�|�B���bf�DB^��e�Y|6_(��~\O5�m��Ϣ��V۳�I�7��z�*Hu���;��]觚C�m�ߝ����_�x�;�ȵ��P*�Br��wӮ���t�����[U�q��t#�N������I@�+�U��(�K'��	�Dv���,��>j(���c���g��-P���u��z�Ů����0YK��n��EK�g+��tҰ��1jcEt}n�{@��BnBE�*�� tu�X��_�=�r�&7�Q���X�8��>%	>7����\�����2�:-j�|�F�`V�!��g�8k� ���F�uEl;o��B�.(�O�H�� ��X��rzy�#3.�%:���%�kW�VNr�-'�]��@�@`��ږ���,S�cO�,<���,��\~.���8���B��1y�"�z�Լ���\o��k*}�����~��}�G3�kl�!�_{.?���r�1s���M���4�%��\���(�1�$�ݏn�89j��\�,_:��Mo❴ʰ2�	�ÿ�����`N,�o��	B�dx'�Q��ޯy��w9:Y�� �<����R}#�Q�S	��}�P�����~眫Ƌ&(K,�鿰:��*,	���r>���?���@s�qu�F��V�9DgU�U���RHt?t�w*o�	��.~���<]��$��V%zWnQJ��ޅ-]3Z��3A>�:lȲʿ��AaՏ�DG]�
�3�[":����	�����i�H"w���a�����d���r��h'ǔ,�+4��0lWբPzZq�dY�Gn��Y�z8��0ag��2�3�I"=��g-�����	�pe��$L�"��/U�5T�Is�q��3�>�������i����Mڕ:ڦ�eؓ��m�b�+���:���m��q�����,��kv{�W��SH9�_����^���뾸����	2�>�G��%>$-h���)ޑ�|����8���q���0�����]�A��je�Q��x�a#�N�yH��9sk&!z2j	D������65��O�Χ�物ی �V��)���FyU%π+Q���lQ�[z��'?x˥����0�!��(5� ΂ٝ'��eӕ2��r-/�z�g�vi�A�m&�5T.9��X�i���{]�h�z5���:���Ka�/H��wq��xoX!��@�� l�1\o�T0)&�_y����6K�l�G聄&�����S���2����D�1�:�������3g%+��J0O�c&�2�2p�EiV<x���
�]~�UT}F�֔��Au���5�5k��&mJ�e9�wv\�H�Me5��֢+���&V�r��X���n�[GF�Y�<"�Ӟ_�r�����ҹ�\G���^<���w��Y�*�C�	�Nl׼���m�Iq�RJ�փ�y=8���L��,6%�35���E�@j���D&��$���4����FnG�h�5k,���j��h������P������>B���_K2��m�J ��2�G��#i��}�V!���	~?�U銀;�`\dz�[�W��.�ܡ�|zA�G���m�R�1+�ޞ�>�Z���Ogp-��T��7�)��Rv�N��l�,�?*�P-f��\�'��ȏ��8�E�|v��-In����~Zѧ�hKq��d��# �D�)tJ�(κ��n��K�4��^��(*�'�oV���&+�3 �ԡ�����K���%� �C>�3����fVh����G�k*���3<���o@|�.��4�w�!�$a��:]\�l�k�D�	.�����"�dg����S�g��*I� Uf��Y��g��{�]]&u��_d��LxG�+*I����+�_��y��{���H��%|��^�m���o��J)��l���/>� I��$�.�����`%���d��f�C_���[mmrD�@
;��a�Q�V��ܓ����~����n���4�v�<����<{��=�NTf�	���Y/.z&tt��!2�^����p���e���Ge�?��m@������!U�ٮ(�C��X����-Bٟ�@�b�y�B!��aUž7�,�����+���蕪RP�H��*eS�#j�2Do���1��v����懌E�� �#��8�h!�7�y4�����&�4(U���@���3���eRI��>�&�-�,*	*O�.y��K�2�E�r}S:�����G���,�qۺ�R#h��P3�ķ6�m.h�+d��~��m��]��{���8иY$����GvAh���"�r%����!
����U��E�u7c[m`�˝����E���b�o��T��C��w�t����j�Ew&M��~����Vc����֔�i���;�t�y0{�S0����X�n���m�G�ҡ^���Hu��'`����$3�L��t>P��˶�&Y��f�NDi���;	�ݚu��D���V�Xƪ���%7~���&1 Iđe�?��A~��=x��Cwm�25��#�r���iC�ׅ�;� e���ݰ�YBfY5iu&ޥh��4�J-VZ��#�C���\�TQì$�F�[l�7�Nm[�4�����������[x��i�Q�.�<S{SW�W��7ob�ՕVf�McZH�p��J���Z��hV����%�[�x��m�0A%�~A��Ah�x��`�0ћ_�L�v�����(��P��6IV���w�Z|�����'�l-i6"GZ/�ǆ);�o��g���F�'o�����IX�7�!�|؟'`;��w���B.�k4�ë#��v�>�$I�?(�����2����ǿ\u�R���x�������^˲E�v/e�P����P.D��3	XtO���d:�u�Zo��:�N,x4c�*�E�Yd��m�ɺt\4L~QE�}}P.gԔ�>%�Dkؙ<c��J=pT+2��&���U�����
�Ij傟靧FT%\8.�����'%���#��?K}Z�����D�Ղt Q�{�jwi.��9�Z���꬝�����l`5�� ���A��޿�i��#h��@k�	�rmRGqQ]��֙lN�^��,�?s4=�����g�~Z:G�4�j�9=�]POe�ו�� p���<bH�' ة7��b�ש���Ίw�@� '�t(�d�3�Y���B�'
�o'Õ�Pl�_��i�<��Қ�Z ��sPFĎ|��Ns�T����'�I~og��e�N�d�/��V�J_9T��"�-���O�l�-��6���nBbV5��,jP��C!&��laa��w1�Jk�����{�
 |�n�v2ʕ�]@�0.t�İ�?W_�K���� ���ߍd���?���ҥ���1�_�ܮs �rL�%Ɖw���8{����di(}v��:�����_"e?�|��H)��,��QQ9�j��Vo��f-'X7�U~�J�D׾ת$(��_&6��V|L�w+ɦ]Dg 7Rw�r�P��	9gv�-�+��!BQ@�Ϩ]�T#�P8������".ws�����?�OC�e�D�ؔ�)�[�y�����$�)��@w"r��fr��~����ܻ6z�[���	l2���IIab*X(덦���.���J�4���)xdB��f���e�������@�2?;a���eG:DH�/'�{�,L��-�P��'�\x��է���g�$k~���)F�h���|�8��̿����*i"D�_����)F)x���A�MY��>�
�@�hɉ��e��04E��ϐ�Hס�x������^Bl/v;<���|;����V��b:��t{��KbF4\;�^J��v�(_0t�Of�p��nDG�����7����;�g�G��q�d��v�ģ��f4Ȩ���<rj��K歪��+�b�<�|��Z����*���=.梑�Hj��!@�.�ј \U�<܀�Yl��mdgٽ�I�uH C6������n7��s�Lh3�>�d�����P���\<�{����������K"�Yb�q�y�r��b]g��l����,���κ=��R7Q� �W=Rc�=f����]��D�F�Ǘg�]w
�����V4�o�2�_�wH#WW�_��b�-�h��]>+֯
�����S�	^�}2|�?�9��O�@$ט$�o���˪�6'�zYr��,��h�t���#�<�����}3�D����ي4v� NK����Ęd.�~��tJ��%���;��"T���Q̕J���炶����e!6�w5^Q!k����<�e]�[&�+�'��>j1�RG�R�h��ȇv@`��"�����_)�Ak��~j�X:KL.��o��#�^�1���u�1d:ե���i1Wk�S��"0�Tv���a�뻑�{�~|6�~��}Dq�mώ���>���%+:��=��Z�da���(|%����V�t�sԯ�
5�ZUq1]���t�?�-V]x�ڡ����/���b�҇l�]w���0 qC����؝��06�Ϣ�V�Q�բԫʝ�J�.j�|ƹ�?B�K�g�Z��l<��� ���T���=���<���|��1$?�~B���
�S���<��-��F[�����G����ײaH��Z|����ԶǮ�&�Smϖ�`�lڍ{?�Y���>W�A㔬d�<��dQ,���J��n��|A�Vx2�$�s_����e1���h�G���Ԓj�˿ fg�=]����n�j��ԡRn�V�/���	�v	#�o?��^���%yk��ʅ�h��a���(G:.8ڗ:�N���S��^��ຒb��F�UHwK�
yE���'���k!��bǎUP��q��
�v�m�g�ȏJ�2 ��4@�&��٪m�蠹H�,n�e�&��$�L�����=+c��e�s�%X�*�`j��є(��f����U�������N�UV�tX/w4�vK�S�"$.�c����6\�J덩�4ZSMc��@V}Y�v�̉���}��Q��H�J���F0H�s���H�3��cdx'�=�m�*^[3GP��N���3�+�؞�a%w[.����kB��������$H]հ��"e�����l�um��{���h
�XPKv���#X�P��*h��#�^Q3PE�j��=G�����$�xg�M
��J��Y0�����e��@�KR_'뱷���������&u�c����f���Z�i,h��vcx�����Oj~Η����Z-#���)!���w%�8�x���zF��x�-�����_h�|��o`��$uQ)
��T�\g+Y',�C��-��0cF�(?0�7�R�+a����޽�1�W�k��y��]���!0h�!�t�M�����T;���t��e3�V���pY���}�8�n�u1
mZ�?Ծ���h�v_tk�U����L�B����7��#��m0_�*�:q�k�_��b����O��2�V��˷�J%�C��J|1A|+��ܷ\�P�p#�b�{#�{N�ř�◬�lA��x����(��y]&�	��mvqΡ���?Dit�aN�9���M�	ύ��{P�᷽eչ��t@o3��RV��|%7�Z�1S�A!���P�I;A�@���)}�f,�qߺbȲ��tBùʻ$Z��I���d@���>�w�����Ēp�a靣��^��W~rxhpC;�6�溰T6=Bc�j� @�i^���Zc�'���~@��eI��1�?'���,A_.NկbJ��!.0
~��yt�^Q*!�u6L*�k?L�� ����g������R6��>q׌����0|L��	1D�1dZ�a�����S)C�f�Y��(���nMFG�_�js�(�[	���z�]-U�a��V��� ��ۑՑ�d��1��b����ƌiF?�~�ұ��b�ꏔ(��\|k�*���C��H�2���{
mҍ���-��	Q�m�$3<E�Zz�U���� ��8*�]0�igY� 䢱җ��F��f��#�d1���.}��t�EA�Vbv��
���Ӿ��az �P�w��M���_���D�j�IS%�<�$NM9�}���u�,̢��J^��B.�:T��S��Q$Z��4��Zj-> $���2�f���(R[�.��a@��(~D��Aq%���O�!e۫�}%q�/�bZ����>Ҷ�|�H d/Q���He}?�VՂ�_�a;�/Ϫ��A��d���1�E\��}H��3��MҐ�u�1k�t�����4n�(1zr�zqŴ����[n&ܡi��.&j
�V\&�mT~�n�7���i0W�Lo���{]��?	 "U�۲��S��Yj����n�O��@�z�R3��k��m�tRv|�N�we�z��� "�T�؝��Z�ݬ3JХ�Õ�� h@n����4eu�M��>�o�ӹ�gӱ�Okh��I_�Aՙ���<��V��$������4�/o�V�	H%�=8J��r՛���N4�	��d�1�6����`��F���>�e-k��tkZ�64�@���,��E�S���k,G)/1F��cV���,-h�j��Qn�XR��&/!GR���f�y���z����k�i:-���@�+dp�3��ٮs���sf���˽I	� a!���1�6ɠ��N��~�u�z�U�y��Tݼ������3�Cv+F�Q�V�v�BcrD�i^��p��A`��<:'̦��`1����x��p�[�^��ܨ}�V�,�	�8C
tJ%����27Tf$RͭgqOXt�TΫc�"�s��].CG��럵9ݲ�{��R�\��r��t\���o�)l��C7~\O��6���9���[���]>j>�
5 ��!
\��[�87lj���������>��wbIX�zу.�*�����&YZ���5ſ�q �s�/A�Ǟ�#��2zT�P�.��
�c�ٰ��W���A����o�:y��M-�,�z&�n��X�G�t��
�A����Zљ�ڵ��ڈ�5����g�n��o����J�Q�f������LU��D��<�/��jib�$x�i��1��`7��Y�MŮ�W�����7Κx�UGe��[E�@�mYCk9ޅ��}����P_.�4@�����7H�kYS/�y�W�I��v���~[��+5��ӟ ��574��:��x�J_�����ra7��pS��P���7֯V�Sn�j�}݌��rT�&�?����W�2�����f�T�+$�1
�Ee�����jc�?]ϖdK#�>Jˑ�)�HZ���?^�V_p��`@�@e1MħC�z�&�
9ۃ'���숳^k�Z/�E���Pa�^;g�BY&�1,�kU��T3o:�@����A�<2���^ltc׳�Ft�0[�����ח���ZM�ek�EuC��-\���ǥ���';L�8��y��~�H��9I��Js��P��@��w�U�e�vEq�|�67Cfr��ȭ�mV����}Q�}��7N:�w�q���T|v,�l�"���Q%Yg~���cC�i�:!�F<�����@���2��R���|��8��={�Mj��~f��<u�v�����&M.�		"=�B��-�L�M#7ZSR�?XBĞ_�:a5�4�ΰ/T���s౅o�=`��֙v-�?��3��h�0/�E�9�J��Fu�jW��-�/,4w�l�=�m���l Q���;J�{Ң@��emT�O�������<�u^]��@���װK�tC�kܛ��k8W��c������9uQ�
�+��6k��Cg��T�CW�Z��E�S�U4z7J̢9�̙������o`'��.��e����K���$-��u�8E������2��0Y���g���jO���Ƕ�v�-z���o�ˎ��8��xq���[�{̻[U�2��?r�9�g0<E�d�{$�M�-m�]�;�__�5��̓���џL�v*l��>�M��.��U�~�KW�dj��vy^'AQ����a9������H�ewP���$bh���"�-%�Q��ޣ�XѦ<I�:��Y�uoP�2,���ds�5f��ƀa��\ɤ�>�v]�o�X�h�Q��A`�{�7�N����Vo<�ݮHT�M�8HU���|��6٤�\�ȃ�!wf���+9�~��\��	K�V={��֦�@W�7��x[D��V�Mp�ODk�T$֬l][>\��6��=�نפ���A-�i�o�5,So�8�t�#T�>l���5Ԋ:�"#&2�Yh!��lZY���K@����5K��_�uw���B�/)�C�k�LŲ�nN8�rY2#/�%<0ؔ�&�ϒ��
�ؼ=w���?�x-7!t_�6,���pf�}OYh�1謀�E<<��sd�.|����e2�k��o��g���SPQ/Q�W�z��8�к����JB�E6��P�|��¥_aM_��n{�:�"Y/Z��:�6�o(��T^1��N4ZTf��޸�@~�o�_+"���i�ͼR����%k�u��AJb�tk_2(���z^�ng��s}u������3C4x|5>T�$�;hdk�T�S*j�yt����w	/^����L,e���/U�x>�T����+��<u�^*o��!|���rm�
^�!�a��Z�(P��ݴn�T<[��ڷ�0��oF��PA�*^o�T��(������JT��������.�'��jmO����w,]�{�l��-�F���/�2�� ��$�3#-�2�_'����3j�*L�,s�K��{��n?G��JNDt�����h���Fu��#�����tte�qNX�
x�|U���h"r����w���/uLew�u��S���M�&�G��Hy"k��nB��+�n����00��[-]��t�=j�C�>��F��x㡶�
H�@��	h��uA��$T���lV!��!��:�c�[D�v��2F��Z����dwfV����Ǻ�ˮ���,Z��ɣF���|%`3�S�bQq�O?ݣ7�ӝWp*�v��ո�̿��A	-�QcFn\��^Z/���4��:��\��%R�k����vuQ��e�����9��RзF�$Z�,�]����Q��p�r;���l�\���@*:�ZS�NíOd�|Q�"OS������_q��E�%������G�r��*���/5��6�ٲ�'r7m��\���	�/��3����e�hOu�
a��g����z�����+P�YP��:&OU��p~�F���Z�5TxUzSR��<P�xXW͈vF�6^YCw���"��q}�W
rq�U='���L��%�
+�-�t;s�m�> _���EG�b	q=����n��)U�"���w��v�l�oJ$t��������U����K��!�,��)��K�|�,�lsy���i<�p�\_� g1�1��9�آOU1�����[����C^�a��ѓ��H�%����-Y#�\�ޏ��_����[�%/���+�y��G����$`2pN �#���A�n����)�H1��(��W9��Ŏ��Ɨ�h���c�J݈���3l��8R�>��y����L��ۑ>���-�����$D�Sٕ4�^*�p�b���x�P)�p1�,8h��l�5�yv��w3�gQ��v>�t����++$ .���m�h�xT8�t��Q*�HXOx�M;� �+�a.�/��AU��_'��C3AdEX����A��YW��Y �Y��מ�<햠z�S�犡�_Pf���rnf<z��}���z���a,�p)����;ۃ���n����t���kݩ2���qn_�9��U,{6���r����nk��R��^�����Kw6����on�v��9ct`aja�6�>�-�\�Yܳ�J���U��Z�N��1�v��	����A�v�`���!�9���FZ���j�5 �E��l�$�1r���(����KN���o���fq����6/[���]g���O��%�S(�!8�����H �l�^ )R�"�M;^�Dc�;(�.y��G�g�?�v�~�7y@IFZ��t���K!�+���>�)�<��qq��>0�^@�{X����.n�y�So�N�ka����%<�.9_�y�`J}pPР'#�Q=�S�ɡ���n�f�b_u\�����
���Bի�Ƹ�1���;8��^�#�c�jOT}Ѯ�k �2&Sׇ.�xN%�s�F�l^���}��O��Ch�S�:�0��;2L7�Ϊ�60d~��!����:�X�q�L��T��pO���!`������t׎�0aJ+V���,}9,5YK�ݥ����b�ڝG��2�M3��
�g��Ԡm�*��o�?z���xK�c�EG�j)��,��C���v��u/)������gO�Ad����Jѡ��̖�5����rIE����5�{,�KN�Gp�d���.����Y����i�����G��3�i�m��S�!�{ꇣe�?3��ϵlY���*�]{��ʈ�}G��N���xgv���z�u	�\�u�W&+d��vI>|4ߒ�>:�l�{�-�뼶ݮF|Nė�s��@C�%z�,Q��E��~Kr���S^�O�ֲ�=��`뮗`��L��_�A��2h��{�(��X)Ar����^��Pi��e��E�FI�V���^J��.i����~��������5s�{�̙�9�2�Vsi�l��Ĭ�H� �/T��r^��Ʒ��C:�ҫ*w�n'u��u�I���E��O�~����*�H-,2�+�����]���{�X����qBRl[U�v�c�bʼ��0�=ѭ�Al�ދ��:������*�[ߟO������ʎ]��"�I=>I]�̴~Z��	�u0�B��~�f�i4����G�ïZ�c���D�B2&	���H���(!�t�!^��ߓ�МK���Vgz��_���;�bE���p8����p�4-�W�RY��:l��y�V��^d��MV�s����c�8l�M��}�����Cz��:�����Ҡ�`�FKT�l���Q������^���F�!�"bNd���U3��N\D8�*Q����wiܴ�i��xwl�J6xc������5��N����s��g�o��퓘�|�^4\k��j�U��e+�� �#���o�l~�K�bz�.��o_~�J�26
<��O|��OǾj�s���4��l'I�W׾���/Q˽��60��>���߲Ɲ���mR����~�5U�b��G9��w|JAӎ<��틒���wv��cgT_�u}�ưo��R<���k�Q��➡{���J1��y��Y{TԖ�˃F�ܠ����ޝ�IWյ��E�;�����1�A�}�S5���:�K�/����No����^���)./1��%`Ta{L�S�8�w�iќ!�\�?��K;UEp��#4����,�f�"�����^V�âr�}���������cN���a@}������˟������Y%�۲'�0��5*�U�Y�%�h$k$e�O��s_�tC�s-��7'��§�w��A7W%P�8��s��0L�ӭ�f��݊����)�? ���h�D��[���ܹ�>4�ͦX�h�[��^�u�	<��=��A��[�QU)�B'��m�D7�}p~���|R_��	��Ζ���?���hly"Nʼ��)�9�/��]e���p
}禢{+c�Q�u#��&��oM|
�'M�`�o'R��~c@3-TJ<V�1oo�/ʾG��z������[E�s�_7�������j��C��!m�_ر��I�+�W��}q��[�7�����(�/��ٚ�b�Ţ]���~��^��%�ɽK7t+�&[Q?砸�D>�<��8L�5-��� WzX��>�E�_�ḙ�nY�O������U��Ӛf�v��輯���M׎��||�VN�'#B��ɬ�d�wj�S*OG���5�V�/x��$�mz_��o��k�<,ԟ�i�k�>ع~�0���J�51�i#�I9�eE�U���z�	��q��n\��>��U����ؖ�v����+Y���	��ߌ^���~��#�쯴|vv�O�; �h�g�jH��+g3�;{��1-�H�{����t2�f�UĊ�j�q�*�6`��H:�U��l&	�^}ĳ��k~W���=/BL�z�=UW��Q�'4��3`����u��v�O�����l��w�(�Ơ�q���,���:�E���y�� SwEm�O�������ɥ3��~���^>�#w��^re�-l��k�7�6�T�n�k����}�M�⋡t���ļڤkV��,�]�x��T��L)l��h�b}��a��W2^����̓��E=˶����?��¿�5X�yX�z�n��Eş�����b�a��dTlz����Ss�W3��ު���'�	�ۘ�XѨ5U�9U�W�D�{����%_���li�[$Vχ��[d��qN�|8���6U�%��������P�ݹW4�7ܛ��.���ʜ�ӌ�d��]N�q�)d��a�z>�(
2�p���w8�Z<�]����z�>�옔� K�VdܼSM�/�h�ƥe_���!�2 �.���?d*f��� ;\v5���mʖ���c]�����O���PUq��ߏt����$;�ӱ�m�R*+���)_}{wsa�p1ʏ1)6�)!އ��O(o��������Ġ"ی!�2�2su5@�B�D�M��ǫ8<}�}�Z-�lۮ���5.�y�܌����c:�7Ҟlˆ��y�������qe_w�x�����č	T9A�fi�I�s��_��R�)h�
�\�]�Qz��X�.v3I<Q<b���o҅Q����ǽ�#eL��N�ԆдR�����_<��=[��.�3Y�]1�;�T3Z����>.�䩔���Hh����߿}����C��)�}����)3�Kw�D��/�����:��A4��u�u��	�7Fҿ<�~]��U[N�6�@��6�4��2��k<������ު@?���q��8��?��_�.~�C3��h��~����.�����˷��L�b��&�"��81�i��5��@�A�e���ھضʩ��<;���?O�����ʿ8�^u�Ѭ��E	��Z;��}VW����g�G�΅��M�*/���.�r�V k��6?\$�k����c,���^
'<n[�:ݞR���`b��s:\툒^����>O���wq+�<�O�C'�d{��n�ց��:����na!�#�+��ܫ��}�:y�w���=o;q(7� ���3:�#.1����v�Ȭ�:R�������	8/L"h�}�F�찜�v�kqS�EU�_<�þ�Pޢ���C�M�ny��T��!���Cn�fw�Bᄠ�6z���8���	��9�ù֡ v�4�"�S��D��]O6ŝ�/+0K��ݾ�K�o-��z� E�Y�U9���4��C�	���=��"'E&)���������\eK웪D��mV�h��������o]rc.��/�=��s눐&�h�IN��9�+�

�9Ҡ����EjP7yaL�
��_0B�/���-f�r�'�-gw�^�Yd�̷��5E�l3��þ��O?{�0j�I�&G�I�˔���$�z ���`��l��>@,j��1�C��N�e��\Z�L6�Y_����Bq������ݖ1<���<X�R�x��GX�--;��_0�=�pZ���I�%�j�sQ�c	����2���lC;O��S�G�m�=~���Vkn	ص����Z֙����U�dndx�����u(2m�%1�|�k�:��~�wbD���6������h������FkI�'Rz����8=�'.9�ؖ^w�9���>��Ǣc�=��ז{ҷV���ND�HI�3�@>H��-�j�~���%׾����'&�d�g��1�e�X��#Q��0/�ʛ��]�t�{53G�f�淽�yf�}��X�6�)������RP(	��h1I�6j��N��V8��0q�bB>6F�]����Ճ�#y��DU1��O�d�,�Wѐ��M�z�I,R^�Cv(7?6;M!+��9U���5��V��;�b��y�9@�K�H,y�	�í5���]�����ka��AQ+~�r?���W�S��D˨��	���&�q]f%ܘ�d��|���=��3���>�1�x�yɞ�ZZ�.7�M�����!�<77u���+�����d��b77��1?��]ՙ���dK�xN�O�����J�wL# H���E���_)��JS �h�a���ګ��eO&�*�A�S��M���zߎV��2�����W���/����DJ<�R"T�VY���vz����Q0 ��r�VY<vV�i�P�C����>�up��͗n�x�h�H��fcfa��^�b'�z�x��xjD�Ā�Xz��϶��@�=> �9��+� ��u� C�&��!��/�.>6��nn������o�M	�H��@h ��0�L�[T!%H �[e�*����7n�c	n�z]�^�e�_D�#��9�5�D�.�/��N��G2ƽ�d1e��\6�%���`C�2��@ߏs�1"{1WS��2#����O͇@��N��^r%	����z�i�R��n��	M�{�h�O�C ��ϓ���`nT��x@��F��	�L>y�/B�^�WӁ�"�v��9��L}1�^B޵xC���9���j�j@X����g��$�Q��ᵲR8>Tf�o-��d�2�~c�H���1*�ּ�Îy��,�΢�?\�{��f}M�hê�G���{�ޝ5BOU�SEA�k���ޔ�
cL�D��� 2��l�V�U��c��T��= �&�i�4t���Be���׫_���d���פ��[�@�q�Ʋ�	�����fH��(�1;�43�G=3�Dߒ��kpJ,v� Q�pOL	0�(�E6��`�,��w<'��="��L�N��E�:=���#�Ǹ�{DD��T��-ݤ[��ӟ���7c�8bB�3�%<��&�Lu_^��L����.k�f����+T#Ô`:ne�b��r�������F�4躣�7�P�}�}8�}e_韪��Ab3�R
]��4�.,��T����P�ig�j�&~��I+��tG`�Ӑ�}ʣVrp9��rW^(��)��0�H�%`|O��ĚE�W��gPc)��= &b�7UFX��v�֒���C��#��Wf449�߁�����~�ވ
5͕xaG�w�W]Э�W��s��c��R*�����B�g<FG
�_�d�;q��jv�d�<��N�n����_��ַ��R��@�x��4H�4N����b� ����m�%�X�pXآĪ���f�^��m�h�k�O����#�� Zu�t��t�>џE�l�_����q���v
�c���>���4 �X��DBcmNr�y���:����xR_A�����iq��j�������Wx =��Mk�}�ݓ�B��">9R�{�>I��(I�W�T��@��б@b�I�%E^�����6���H4�@C�	n����<؟';F�X��^��}H��!�s}���r�A��������x�/�r�p6��V�����L�県/�%�W���7aor��VM�_��"����Ӈ�F��Ԍz��J�}� M'A
;��3h2}�/�~{�,����SN�뇀����tG�.�/���#0T���-o6���+�@!�$��-�ǁ��7�Ik<�o[�m+����s}x��{�A�?=�=b���ƍ��m�Av�}�0�Òp-��!Y�R��k����a�����K����k���I�#FL�4��l������vFT���T�}� o�E��BrlE�`,�<6����C�ܞx��b �e���O 0��m�xԂ�<�l���?�%m�i����L%5�Ф��D/;v~>���Ɋs�l�&���u~�&�����d�=xN��HM"�DE��a�ee�G�����%���o�A,b8���;kb-�=�ef�wn�BvGn�N,��� x��>�x��K\o>��q�t�n�L�c0�[a����c9(b!��)���J��*�?0|�'nnx�sX����.7������qv$ P0�d:�	 ��_RX�Hx�����@�	$t
��^�e?g��!�Of���^�d*t��X]�b+p��Ԝ_FG��g�C�T��ё���2���ު�S�H��IL�hڎ���,�G͝<�n�^eH��7���,��ZC~���γF��&�в�4Lg�M�_�B��Y5�i���l�w��sg��l�j�fa�O�+��/4'>�Eٖ��֡ںУ�z���u��mA�|J��7�f��
52/|6>@3�p��"fR4���$�@�^�Bg�.).SR�B�YU]Lׄ(�8��f�$?t��R���#K��g��4e����z��Nr��d�l�)�> -�x�(�z��T	��v��%3�8 ��)M':�使*-���i�a�j�h�Ԝ[�`P�bȔ�:_$�vW�,u-�?����C���	�#����vv%�1~��Q��/�b�$�=HR�'�������R�lN�;` � \׷�̝ڹ��5�l��<�Jn[���z��f�/�0@�M�!/��l4�b�)�k��L���D*�z ���wUc��l���kX8�Ŵ<����e�`d�D���wU���Օ����@����l�c�ӥ���M�M3<�P�ߎO���g>=:-�a���Z�rf�&�W+[�4����G�i�7V~D^��D΄�^��6�޹W�b{1_�o�C�}~D�P�Uy�F�(��*9�����<z\><:_Q�v)��q(r�w�r}Q����YiY@ȉcJh3a��]�B�勝���7%k/�bL�bSt&��S�����`�>�	t�E�a�r��}�"��,2"�T�i����ڒ��H,}ڔ�JY�DɥD��������ts��E�Ŕ��`��z�dcęɆ�rB�UYO֦��N�~��q#��S�S����㋹)~^��R��wv\��M�73��U����̙/��^<�K*џ��!��5�o��>5 ���+0�� Xe}����Ƙ&���7������$���nxs��h�\�!�A(A>`J,���XF�p�'���*V+C���G-�N��2�$�.=����tHP'46w�d'�<&�K�oc���E��̒��,~iO�ҫf��*�ĺh��XXLQ@�c�Vz�-�3�#�?o�xid^��qO���
�#|�y�b�f?�!�8H�	Y���87ʗ�w�A�8h����ͥt#��0r{C�\{�T�j�u$�c�K���0�߹wٟV&q��?�Z39ɂͿZ�W��	��DO�NC�����GӉ���(}�����[.^-�&�v�/�������Z����<-/����5���hz����mx�-���gfA9���xO򎱩�j�c��+���f[�q������мI`���vzԮ�,�K�Yn(w���u�8cja�#rx�Fb�qa�^�I�����|�R��
��8 mQ9�C=��XzU�B��N?��L�8�663(�l�;��xv龷���~�lOTs>���j���̚VAo���C��i�Ɠ�N��iӧ��rg��,������3�2wt��^r���Kd�����gA�������k����K"��Mw��l����q�>�^�z4� �==�0��0o�T���C� p�ۘ���~�%no�?�`ke�6���`WL��8π{�3>�^7�iDc����s:XZ�{ϔ4�{/?G��$=*�~��o�|��+-<�4����x>�*������� 	�$�Rz!���+	�yֹ������o���+��f?��M��~[��u����Hx""x�~*��q!%�'k[{y��/k�3Y5�BpO����E�6�tM�0�^�=ϱ�7��(5j�1Լ�j�%���
C���G3�T��y��8�q�;��^;Ld�X���@-˟����d�xCj��So<H?!�2�&���E��z�J�uo�BDT���(�6�ِ�(呎{g��Zl��ӥ������X~��_ֆ��tK9b�H�5�l[FF�g�H�ӈ{��!��y��5��$�ﲈ�W |�δ��܌ˮl�'MMT��df�TD5�����Oj�C7V�� � ���0��3T���r��̀?с Ƭ�p1��B{A������H=~J}���e�/kE3!��nD�du�>�͊����Q����zd�=��h6����l"����E�����|e�,)5��J3��_�-<h�9�O6g*�j�/��&�ǻ���Lۡ%Tآ}Z뎩m�,�c�LM+���OҰ�^;�h���>1�X'!g��)V1�_�1`�x��«�-ue~�d��9AH�[go}��; �r�]�E����E9>��F���-0������W�����ˡ��Uh����M����-�rR�C?c��RN�5�ĕr���fX�R�ڿN�5b�#J�y̗la"((7�@C+"E��x
�{�:ݔӍ	��?��8��X��[�׍C�g9*���!�5�A�����2j�׬HH\��)��s/EI�HW~�~�C�6�VLW[��y�XABS�r����ުnƭ �ڜ!)d���t�8^��634����:;���'�259����;��)Żh2�\;�}���Ԋ�-N7&�����7@"xV	��i�a�w.;����s�6Pa37��1ø �a���R)�� W-H��]�C�膾�/b�1��=�J�æM�aDl&�X�����M�'�|�v����5��ϧ���Ҕb���p=`놡��:�	2������//"�}���%��NNi+)��u�� ����,-�I_w��y���o�]���,��]�#�\헔V�@�~���e^��k���L)щ9S���ߵ5� Y��1�����z�X��� [0�L�V��ʈ c���^m��oԼ��1P�"�G�$3��Y�S�]6��[�e���)D����t�{l��0�Z=<;���ODz��xE8����ɦ����2v��Ks�Deca(�Ki��ɔE��3j��?�_�h|T!Ik�+P�w'C�'�(�������HB���P��{��eo�v���f� CK{��O�^�,bhQ"����4"�P1�Qک�v�%+�H�9GQL��r#��*{Z��aq�B�1����#��ܗ�h��������Ӭ�;g 1��>o��s��m��B��.����x�~d�\/�$��ds���u�~�K3��%��5%��ƛ�2��Ĝ|�v��fE���iI�?��Ήx��v�C4I&c�o!���Y���{�!L�Xx�#�pE�k��
�1��ί1����z<�zUn���')3���$θ?U�� 2��J7��1�@�#��$6`�;����?p��e�/��D����u��;�|Ē��>z:��B���8�LVP<�joI��r5RE,l1��!m���qW�U΂pS(^j}�F51��t�����.���ۿ
F��$3�աN=p���r�v���V5�dE�&яx-�Q�-�R���c'Q�$��=f�C���s�|Z��ը��R����KnI��!�Zi^^���ރ	���	`5uG� a�?�Ğ�p򜄟�>-��Q���eJ�����J��Ф���!]�u=;�"����s��b�o�۵e��@^,9�X��d��:����%���M������2�M*�����/W�s��LXڍZ���_���/�F��h��<�m�xV�V��U�~�L��D���.����*;&<�}"�;�v�V����IËb��¿ߕ�.��P��WQ�����oM�~�.r���㯹C�9���Jީ���`D�~�;iQ������|�ܦ���f2_U��6w8c8N$��AV;{<���_��vf�!��Ĝ��h���I�'�(�t���0)Z0�08t��KX���R��z�}�t�v:异fcT�[��L��c�v�X����B䇀�f[E5.}�s(b�!/T᥀��N$��儣��~�"��U�ջ��;_�.~���8
��ʌy����=�}q�q�Sڞ�k7�Aa��ޭ��
u�]<1�f6����;�O��a<
܈/� h�{�m���O��c2|آp׊Ex{�Ac_�מ;N�@��v��?8G L��V���T�a!rk
rA�Ƣ�l�L��G���'�������yY�?L��q�w �F:"A�`�͞X���o�s�� ��[K��B1z�}'����s����ӈ^��������*�"��Ryg��\g�eQ�Å��r!oגi�r���t��)�PAP��x���(�Sc����\���~6Ԛ�t�M�e��C?�Xem�?�=xv~I���к��f#�yay4
$�h�^J���uh�L���*u�
h�{�K��cw���0Vf�v�����q���G��j�@&�̼�}�Z��_��~2����83|�Xs��u䘩z���G	b `����\�$|	���D¼�BM�c�^�J����]t�L��p�q���m��#�M��KB��.�\Z������M״����d��|�L岆�G�ח7��Yuޟ8��5���t�E��$fᖟO����I�D"ux�X/"���f�:
�D`EPA��K�NО`G����Rt �j<jip�)Q�cX��t�9*w������OG�'�4q2�UJ4'W�B��b�<L;t�
�)�W��X���!��a��PVaNܽ��եVÂ����@����N��a~���Ǒ�cF;�<0=?!�)YF^���pt�[Ta �HCÙq�P�s���g���a�d+A���'�A�}�E�K՘l�]��;o�Q-0�Ϲ�{ׯ������iu!)��h�˂�d�b�W��>lvUh�I�/���5��̠e�l�W�Fxt=���r�g܈�<k.�+ )x��E���w�>m�¼�"	%�!�At!��5S)::��m���������7��-Ĭ�n��E��t����^̶2L�_
q�Y��kmSa`+uT����}�s�� Ǫ3����c�2��̭�1���B_'�'{�U&�g���9ͻ�{�;8\��<�8��)Y�H��8�U��	?�~ŰV�'����3LZ���j�VFG�����Rz��kՃ�3R��XQ�w�g���!iK�?��������!��:� ��>m��!E���Lsq�Uy���ճ٥����g�4�L��#nL��%�@����Nr��_�[�@��+ҁ��萣m�_�����D�\������0N�&�헆��%��?�i,��5��>��^���*"?
WW�����϶��gY��K���_E�	�'zڛ=�Ji����eeM�]��F�8>�� �
J(�R�M�V�n�S��~�S�-�,p$�g/����}'�27>G��-Q����/x�b:�cy!dj��3��D�e[� qy>��J�{i?�[��+$@���*h�#,^�� �{��8�����;΍9�#Q�?p�p�DѵtŸ�*��-2���AJ��8vuZcv^��V�4��Z��<By��#䛰k��'S��5�`��*ײfN+h�+!+�o��b�F	8�H�H�M8P��ll�Z�7��j��8�8��i$*�7���\X��f�m&�����Kp�f�s����4D��]��&a�n"i9�%;7����; ��:�1x×B}��B�M�_�It�M�.�8"�Q��&Z���!��;�Z��d����?�&���N�s��f�J!7�za0zu��,~
�I��U%�~7k���㻎t�q>ʩ��H9dLrV��>â� K2vA�"�vC��q�E��%#Ƥj2�/0��r_���~϶=��Z���9뱕9 ����{�&�\ɉ'���x�9�/Q���}?z2䥶�׸9[����Α�Z�_�ޠw׀�-�F߽��8*=,�Bc��J�����w�1�c5�fX����Z��)}?�}/c�2m+���{�ͳ�#`�G�Y�����	�ڷBT���2 ��j���0��C�jWtc�<���q�0�:��8ʐD��<#�a;�]��I��Z�oGn\���/�4ω�PڰIz6��H��;
�?A�д_�)��ۦ��Ugy(u�x"j]�B�k��z��WM-�>ې����m{��Dc;÷p�I590�T�԰����v�h�g\���2J1T�r��M��{�o^��$��ɽ?���OARS.F�ϡk�z[�_����!�6p��ƠK���1�h�	������f�>%0u�	��߽(�I����7�ǔ��q�`	aQ�P�tH���n^0�%�`S��_w�h�ۅ��ܖ�S�y>�lO��/��g���ci+��#�����y����#S��4[rS�ށj�$񲇋�7{���/�Ӂ?�Y�Cm$���x�($�f{?�e�b S��/�>ei8L�2fe�gn����iX]��IY�_?�����0"��/��r樻W�r�L'm��V8`�.N�������9���ٴ�r�S6o<���I5a��P���/�C�a�h�M0��)HpGY�J?�w���]�B���N�l+�����	j2h����0\��״���n��j�iR�o��Waޙ�mg�6��?Y�����U�ɑ�ixs����%T��{Rݘ[<c�� ���=ߔ)a�?	EN�#�" ����6��V��q�V7-�?VW/l�!��z���w�J�+Q��	��#׶��C\�[��_��"�ߖ���{�������^�u�����7���&NF��bg��;��X�� e;�d=*2��� Փ�%9��≇�n<I�gNF��>�>�I�;�T�������(W�����6��e�� 7�)�+)�)N���#�i鴯VX�|�O����#�#���f�us_K�q���G��*凞'-���ʿ���X���g^>�ۊ�NA7
*.[d)狙zk���Z$5Z�}�į-7F�p=�[>190���eN����b[UqY��Q�,Д�Mn��?��!�z�<����	]@� �T�*�\y���9ǯ�]n&�v��$�]�c��A�i{M9�iD-��3~��R���C745W
u�(9�Ɗ���Tu;���|X�\,�:U���D���[7�M�'�7�|&T�@Df4[ژN�T?ks����D~ 2�&�t~��&vo�?8v��	Z���=�Qm�~���?�Lc�i_������6
1�~5M&�o���v�k�9u�D�y�v��p��Ld~�����������~�H��U5�ʠ)�W<ri���H(���g�Ai/���}���JD���=wz���WH�a'��s�2U@�R����X*1�׉q�ΨF�ï��ь����,�9�	'B�wh�A�UE{���1سE�IC� 2Q0�;���g���"�̓o, ��rEFiM�K�-b�(�M͐�Ӥj�cG��ˡE�B�Nn��i�XIQ�D�^�8T~�tk}�*�Vbܽ	ʶڈſ���l�,�W3�����(0K�A�Vɚ�b����r	�օş�UΌc�Kl OO��?W�kʶ��F��SUez��O{	�i~zY�"���m�F�|	v	����`B&k�Ϲ�0.���e���>��X�vH���Z������er�l�`��0�p��6p�K�ĥ�7�g?���ܞ��8C�YQ����g?dG��%�F�q]�2�%�Dز�$XE7L-���D��|��Ti�Xg*�"�=��_iZi!?���q��y�?��J}?̂ć�Nݣ����-���Ԍm&+(�T�T������RQ����^䧪gR�<�^�	Rh�A����W�#��f%�N;O)QK�Y���뫜I�1P!,}�6�
J�
_H,�sr��_p��(zw�a��ą�U~�q&�`{�l3RO��������S���w���I��Ҝ�O��Z�j�
wg�i܋2�0.$G����01��>�R��b&�{�m#�f�[���Q��D��O��Du�u�ϟ�s��R�N�m۽��pv�m;�3�3���;��2��O�����|~u�BW?l�yɳd'	eib1�;F)����\���\a	&�W���k��N�v����9B-�5��+]̀�.�{��x�.�]�j��?li�Um`�TkKrQD~�c^x��u��L*n����Ad�& ���=Q $��D%���(�E��Ⴧ�{�w��k&%�&���b򍓡d����՚�@�F���$�h"?�aY���U��,r����?����¢J�����:�����6��UF--U��}(�=���`��*O�z�m��)��X�^2|�M���^���$#b�~�n��(������e�;��<V�k�)҈�C	�n6�)ÏЂO�ƩP��W��5�iN�7=c��y�>�c׽�e�UPm�7�c^h�����Mr1E~`Wm��T����� �2_{9n'd���t&�k�d�B�*���I�����ʬ][B�r8۶�}u1?P
�ɶ�&=��������Ђ����R���ey��üzۃ1�\��������>�x��-r���*�`���J�t�w�N��b�,ra{M�KI��w�ך	��Yo��jVo7PcY���*H��I��L��sq�����yS�)?&�ۛ������oom�(�*))��<U��������3�o�p���UV�9�b�%���_̾�M�s�I�*��
�c�����p���>�D�~�਴C=8�=��[����L���c�端kk�*2�>�055=X3�U%��Iz���I�����̣m0���"r���C,5u>R+�O��,#g����_���_�Ԛ_n�YG+?K:u�5�41j�O^G��,�j��qzz�C��ɟ��"�@�`���7;���/����{[����}9��pɸ�}�@܊
VG+}kY�R`�I)���ӵW� ���p5��`Y�F7�^�����x�H��ZN�M��˃'w���߀�>z�ɽ&�H��0u0�AY�xR�;r�c�]�f��^ǽ�6��3�>R�tG{������ߌi�����*�//ǵ�朊]Ǎ`K@���n��e�z][[;2���Ǝ��j@N� �̵$����ZV�MF�f�P�~Y|����	>Zxi7>�&��o�ԓ��Ґ�)��~�^T��Ĉ����/{'�tCm�ǚ{S�]���ES��wx9�4GX0SΟk��?ow/��ۣN1���J|��|�0y��m�������=��B�"O��]j���8�;�K�G/�	ń΁�x�Vf�d�)��K�߭Ś7�v��˾U:~�U��[�cI�s�/�_����ma�����L�~�|�onM��]�ï��m���)����ü�wФX,V�~aѥ�T�xO⢸Gs,A�=�W�l��.9�B����9�������;iϲ����n?����0�5#Q��C/�C�$j"�&����U�,�?�`m�/���8뙟�ğ��ΚR.�v9U�f���Ӟ�Ԟ\���:M�����:.g�40=��:=�:h0���x�8���z��}�b5`����p�RP���9�Y�A�9h��+��Q"*�)�9mA��Ѹ�;�]�-���ѓ�vȑ���� �R{y��s:�J�J�@�Ӫ��m�a���y�L��XRς����u,G��썓�6?�־󏩩����H^�����F��ތo�6�s��[܃���KR��m?P�.T��Z5�W�ǋ־�g��G�%��f��4}������v�4vs%l՘Z,I�]	�.[�˺�o���b��	���l�G�@X���鿟�'�*�[��J� �ul��J�xR���	�6�b��8�矎�?���ͭ�G���Bz���-3mf��/�?p��9��F>߱m	�Ѹ��E{�G�>^=X�΂�\_��=����%�7|�h�$��������6�֚��^��.甌�Q�e���1y�Ӭ߱S̘.g����/ �Q���Gӽ��'�}�m��G18�;D�b\8WL��n�X(C���?3o.{�3�]�,��?w�`���䲭x6��߫��
���L��h7�9d�=q����ۤ�U��4Mh�
��=XqFi+-�\2�wU%��]�����UC5C����|�n���w^3>�"��?�����(n��Wem��J�i���j���f؅|��;��"�Ƴ���T��*��J�ߕ�Kv_��1�B@HI9��l�����=������5K�DX���C�-9�5���(~rz���x�}�oQC�	�1�9
���Ts��p����4~��V0�.5��gs(�*�U�l&��Jsp'۲�ٯ�����2�ք�5Y��,�}�`6���w�/s��?5��N�J��\=H� JC�"���1ɶ��k����&1�B�Rښ�p���12/M���z`�ژ����}��&L�1`���p�EA�4_/����<�;[X�LN�9&�$f����`ɟW9�1����^Z]ר$#�依Z��$a��M����f�R�].�����	��J���3�6Z�.QZc5<�oAm�^��_̐�ӱTܡ�6��0�	",�LT��ިSk���'[��t�m���J�w�	K�D��~�}����b8��<g�`�����(���k�i=f��f��ge�e��sooG�B$�s>އPٍ*�]�>'lK���v���5�N�>=��U��f�r�Z�P�HE{l?Mulݶ"h��`���W�rK%�d;p�*h��]��c��>���� �Z��F�!�����)8l�s�c��zM���.�Ss���s7����Z���s7{H5m�hY��2�Qt�#YMV��Y5����!��CJ����N��K��*04�e��e��2�W�1}K������#�/��]O���ı)�s��,R�|������mq"�ŭ����7gH}� ���\������Ƽ�|U����åa��G]2�z��yS��+��8���<��T��ȱ�����I�s*�y��%��{�~����|za6d��?�Ř�~wa�!�3aH.����㨿G��'8���EI�`�2�tM�}�J�ZG��?u]}8�{?�ǩ	�y	��^bޮ�lu�p�[I�!E�Q����UrD�gΜl��y��E�$S��ቱ�D�"�����빮���������~���}�׵̓�\]sGt�Y}�ܻ���s}}};�@𴯏>(N���]l�E�f��74���_��T����&R;��v"wL �������}��ir�T��#�[�}ʶz��;���9���g_~��� TOhU%����`+`"��q�H{N,q��˺	��b���1��7�"�Z\�f���1�ͼ�_f���]2ƮQ|���E��8+F�Y
�GE��x��Ր��^��O�����x|���2���;	aaaa.����jO�)
_��!�9u���X��L�����g��"Ƽ�&p�����e�|Z����7�x�uX�G`xJ}��:�4�J̭i~cQL��g�ǟ��Bd�i�.��n�?��
�e=�@�s��=��nO��g��s�I��Za$���n��O\xt�.��g��>�Aa!�K�Z�T�ȃ�J�Ƣ菕2ox������6??o�΃�Y���E�m]��p��0N�&G��|���=�F1T��[�D~�>�A�32z���A tt��'��2�&��,������!�	��jX[mm�j�=�z{����%BWi:���@rZ�6i�ag�P-tr~ܐ���^��>�n���d��|J�^����m���IM"Mۏ�(O������ᱝ�n�P!C�Z����_�e`&�V�Z�$R��5���s�x�(�Z�$�/I:�s�rgV�8��:@6��,��q���p�J�cRs�.2��A�ԉb�(cP�d�i�
�(bR��W!�X
��d�n�@�ť$>�
��!��B�d��������B��9��~ֵ�^��D�:�O^y$K\�+�jA8�<��q������<7�o�p�#�PX�x3Q�t��=�f�tNA)	�P;[d���{z��c�.��#��N`�7�8l���Zzr��A#�'F���4kX7E��/�Y*���-Th�x������,��g?�rQD�uE#v�i���%#��a�"��6Y���f�����C�p�)v�P�E�_PD�b�@�@)V| x������y��H�wA|����b�n�YY�H�A�U�N�0PD:�z;�Ig���M(����1Y&#h�$m�=7�|(HG�Q� d�Ce�A��Q�u@�)I�Ǒ����B�M穁"w)��啒���o�9��8��^�<��vK��*���@Q�]WP�1�c�1�"����9�%]��z�����i����:\�w(L���u5bǃӊ�9�t�1�BG�1��%h�t)��=�n�����6�gW�T �0�������w��HgO��a��Z���C%=Axr@͔�)�X0���%~�|�R�h!�����5s�C1�j���u���u(�F�Ja�Yv��"��s��������)�.�!��;���q���r1�]���R��ǩ�W���~¤��	>�+��^�]��~R,O�%�@��"���͑�฻�W�x�aM E��2b���K�;^XJ�P0���k{�k#V\aWղ���z���J�6������Ƙ�[~���W��]UQ{R�_�P�$I���%���(���c�a�{+|�<��d4��ԓ^�d�k�ys��m[[r�?�g������P��vWd=�nr�R��e�q��+~��%^��q��q!�B�̅ ��8k"�m�Դ2G�D�c��]ϙ�\�}������� bVu8��t��|�P\�pao����W�F��j�h�%#wX� l3���E������C��zg�y�2^&���Gͦ7S�CBB�A�v![��.e@_P��M}MI�u�1��'�x���xa'XT{V(������,2Tdם��eN��pifvxyR�����!I�d��j�H����͒����O�^n[���`�:ֻ�&��
&���TuE��W}`z�p!���}~�9��o�Hq�Q����k+�<�oH����;��#m��@�Tj�>�<׺���֣����ۼ2��2�(���6��w�#r��6����Ԙ��Fi����O[5�iT�e���U�k_ e{�Gd�8�2�iF�h������,)k1�������K`+eڷc��B���(��l�q�{��PK   �2>Z Nu
6  �     jsons/user_defined.json�X]o�6�+��6��}ɼqP[���CPH2�jp$O�[A�{/��Fѡ�7K"�!�=��O��q粋�0�����M�6�2�����Z�@s�3|3J?t�.�|zy�.�ܫ��?��5�8�*���ql�^���[�@/�����Y��2]VI�D����%e@��T�,)HyZ��U����5���4>W�,�Z��ԊYJI
����X!]�����5U�'9��r5%�,��(F�p�P)�嵖@�ˤ������6��[���X�'�_1	oۺ�.����j�ݶx�춘���\(��NN��w_�7&r�����D����}�����cE��nh<��f�r�rc ؒ	.r��4~��Om���q�K��E������y9������e�3��b;|���� �Y�0 �Ms�R�t���Q" � �60AET���
�h�"�Ab �>AD DXm̩�gɄ^Z[:�\Gl��ՠ�0�� q����r�BY:����BI{=(+��=�8�X�i�M��s�\b���5rF��\������9uX�(B(jl�:�Tr��[�uy�Jg�j�[�¦���=Y�s&S>�N� ����֩ ��L�SU
��w��,~��r;77��d \f T�ظ�J��8����(���t�x���327�(M'Q��|�xf��߲t��l��(�Ρx�桌�_2�X�Y}(b���'���L}Ck�>SL'7�s�����}*�H��Xc�o���Kӣ%y�W}�s������]׺v�~1E̯��������ׅ~���͎�cD��"��5)�6����X��2�D�4PI����ݔ�j
G��0R�Ơ��P�M�STqE��@JM�T�!VZ[�]�����A��f��Lgx�+��"�`�69^�;o�֗�3<&��AC��$u�AC�ᇄ�3Ï�LL���� �����Gr,�]�$a�J�PU�D
��5�򿔤�Ve�7�_5�>�kw��^ጘ$�w�f�(��_*T3�5p��3�{��!�_����SpH�֊O�)�r�w�_PK
   �2>Z󁁣d  ��                   cirkitFile.jsonPK
   �S;Z�%�W�  ��  /             �  images/538bc4a9-05ab-4361-a8c5-43654019cbf3.jpgPK
   U^'Z�!�� �� /             5�  images/a017e9db-93ae-45d1-af88-7a97bedfe2ef.pngPK
   3)ZZR�yHS �Z /             k} images/cb4aaf6b-8f50-4b44-a327-f08934ea50d0.pngPK
   �2>Z Nu
6  �                � jsons/user_defined.jsonPK      �  k�   