PK   lV9Z���  z    cirkitFile.json�]K��6��+�kQ���nc�l��vlox� 	���jU*�=���P*E
T��zǮ��@�!��x�>[�_��Z���/~��X-g�T��>�u��u%7����n���i�>�n����_T�O��_n�D�x-dUS�B(�RKQx-m-�6V�;2�}�����).;�e��"d?��6^Ѧ�E�]�ʋ�IK
�0�pA\���qG+&VRnJeSj��օ�TV��B�*��k�k�J4��ʕĈ�1�,��p�WEU�JІ�V�T�A�F0�1-F���De�c;����"G7Eo*���#�*d~�̏�E�!��hb��T�\�UKG�wA�	#eȭ��4��V�c\2��j��ډ�S"i�K�eȭ�(x�JoS��ȪSb����u��Bx�
�)�a�)ʭa�)r��Դ晵MY5E�G
�.��U��U]�P��$��T5N`c��Zm1U�Z͑z���5���lDԜR��!��:��CQuJ!���5���	[� �ơ�`�ơ�b�N�1�Cu�k�C��0u�kk=c��E�P*�-��lA+�-�DCl
� ##5q *D�5�k�ț�� �(%c��4�0�1���|�6��\�:�_8͙�@U�?"�p��p�t�64�,UUT��2�`-I�B �S��g��`0����lDͩ6���T�A�SmFiOP�(9��Ѝ�ɔ��:�eO���yQ�L����bl��&B(�k��:5&�Q&��H�d���#n�Z fH"�N�*�D���~��Zݯ�����_I���h�RX�Rx�RD,�i�5������k����u����4|i�R���<�y Lu�b��A1˃b֢��8�1�lQl�lL1-�)�r�U�Z�����l�b��ӢX9�T�)f�b]�SL�bKkRa���A1?���K:�7tyf\�Е�qiCM��� 2�/��q�A��q]&�h�>C)���/���+Nh�w�hvuЈ���������/���	�������A���v����Au�&4斁��_�)ACb�@CT����w��O^N��ُ� ���m<6���O���GX�,��,��,��,��,��,��,��<���<�y�K����0̓`��4�i�<(fyP�2��<(fyP���A1˃b��,�Y�<(�'Q��K���������K9�/� ������K9�/� �����,�R��r/� ���-X��`�������X�4@���R�|)'e��K9)#p�_JWF_n�?�l���-�_g����>/�����>���n��[�k��ݾ˾ǧ����ق��z��
�WeU�,�������S5����B3LMiaIm�m�MY+*8�f����2U3��VF��$>�KRVD� �RJ+�(Q5T͘ަ�@��K�Q�%j��: 4�15�֣153����#����$-*������j~�6I���W�[���n�l6̑C������sQ�MۈOFEz��7a���I�A��������5)Em�K��;9��H�İ05'N����b�9�����a�@��LS�}U�PFh9�S��p�5�HR��xՠ�����_,Q3�l?�����N��9=q���fkP��Q)�(�
cBx��)l�+�8�J�1@U�j��:�����gh30L�6��`��8�σ[�����I�����JE���J0ggꦐ��Fۦ�JO[�ܘF�&̳L��)��W�Sf�C�ɚ��+g0P0_O��� ��xC|iHvs|E����7�f̨Jb��ڤw�Y|iivt�/i��.	�𼈼��V����-�c���W[U�+G1�\\e�k�x�Kͣ\b�� r��l ���� ��G��j4��4���4����*��J5���(Y��2��eV��;����pQ"��K�g��W��&���o��ާ*���X�a��������O�2{2��݂��.���.�#�m���n�J�><��"��%v�`���T�TB��S] >�3p���l-��(�^ӌg�,p15C�zF)�1��A�g�5����B�-p���!��[��7��%6��{ ��od$\��S��Ev��p�M�x���8H�@�O�dX��
P�؄�g ��o�<_�b1�C�?o�nZ/��2v�(R�ܓsXh�-��\b�jZ�&��C�H�+�z2z^N4����9Ax~�w��+�S\J�'� ��gx�',b�F���n~�Q^���\«�|���6�(�ez���8�(�8�q6�z���3gR��s��Zȃx��?��g³���� g�C!�UE-?��ܺ~Z,�;�WϏ��W�5�͇;`(2?C�����Hr����By������N�þ��i�ł�V,\)���1TX��8�
���@�X$2,�'z��mP����fi��=�0[��l�j)�H�P�R��f( �;�4(/������=���;��ک}���S08��|�56���X߁_��a���w!`}~ "cqG��&'�;����j���;�k0����1��i�~h�W\j����Ч'z�a� G�þ�	k,�U�^i�Ǝ���)2v���T�;�0Q�����s��X$D	~�"cg%�/Z���c)���H�mv�ny��q�P|GU�o�8]G��yZ;� ��Ѯ״��Fr�i�@cs�Ǐ�(b�Ǌ��V's����,��1�W�� �Ԑ��bG���_2���<�T�4w��U�:�F�Q�.PV�KQѲ`�sa�r��0Xg�:�4��Qf�& ��asC&�$uP�¨�y�ބ:��Ѭ0�g�&Vp�`��aaJq��GFAԴ�UU�@[o)!s���Ft����Ha�=m���o���6d0�o��bN��y3+`�$j�ˠ�i��Qk���}@�c�b�_�s���0�3�NFm+��$�v��U�n:���+��qn.�
�0����0���>��e^�و�*��/p�&�0�������>�qn.r���8��E��:tfзj#����Z�b�n⣆����Vi�Ǣ�����%��^
�%�a��%�a��%�A}��+��ʆ��+�mV�vij�M>g��ll�ƆIϵ�L������?Bϻ���r�T��:^�٬�������h�h�u��i�\Yp�o����w* ���O�w���7���D�:n���Mto�a�z���·>���e�_T��q�^,
-Y�O�;���~q�O��om��^}Z.B%��Ǐ��o�߆rg����!�ѯ\<.�{��m���i����ۄ����O��6O�x�i��.Y���f��VV���b��]��ky#�\�?tg��m�x]J�[-%)� U�+S����Z����q��6(�r3[�A^n����!�T-�ս�I�]!��Fȇ�ȭ�|�n�즈n
��N
�����Kƻ)��B:)�vR�T�0������)���m'��n���n
聆Nʶq��u>T7EvSx7�uSH'e�����ϋ���S�X��׏[I�9����#��߿/���~c��[���O���PTZ�,���&�!Ȓp����u$u�]�`b�6�ta\-�%��m����$(X�r���v�D����	sD��_��d�q�N�E�9!AW����0��o�+-�b����yȂ�<7AQg[�յ;R k�Y��]�X���C8�.������WA%�������5���/�-맘'�$;6�Ϣ����o��sA��J]����B�<`˹Bk.�5��{DW}P�V4 ��=��PњGZ�0J���{`B�~
\����Ebo��������xXݻ�b�[���O��;��J�F���+��5���o����?��?��n3nJW���z�������w�za�O���6��x�_��yp�aˏU�L������4�/�����Y-7o��GK�'�e�diɒ:�}�z
�a�����1�6��kB�	޹PZU,��3M�іٸ|&��YHÔ(Y�x���FxË0�8'�V�4���xz4_l4��a��ϡ���C�E?��m\���n,Rƅ�Thi�{����3��I�T�?�)���Ӡ�ޛ��u���3���
�5���U0���TT\�&��t��;<dF_�mto`T�6vS���}h2'J2Ev�;���?o�)(�J~89��C�Ra�U{C��9�Z
����lXa���/�RD{��� ��8s[�!>�[{�����#ߗ���~��\\PM7�9��_�܈�B�=� �+�}�#MU��%а���Ԕ�A�؁� m��Cb����}A�^���so���Rp��0i"ߞ1��s|M���s˞��!������7X�kR*��JF�6��&L�J��2�	SR`-A��ȯ�+��"��?�SƯ:5�#��*���sFy0w��ez$�v>�Ű2f�S�<��`o�g+�c�+�r�;��������'V��U�f�-c�2��6���)ʤ��ù��`�ju��7����PU,L�H��`p�r�X�#����k���r�kƎ,�>'�t��&Jq$��h���-t���^����/�2.2�tD.�n/D~y��~
��Iv=�TH�N��<�W�N�$n���m�`7���f�TrNä�g��8�F����f�a�7c,�~*^�~��[$�cb���1N�� �o�5ĳU����o���~X�����?�s�q����p���~v�>�qо�ݼح�Y���n�^} �-�/�Ѣ`�%ڢ���ۜ���������"�n�-��������7�1�m;�=�_o���nw���;FH�!�7G�x��̲אm�<��	5��&�=/�v��J�d���}	0F vd�*����u�����"<*�`w�zL ��8ʭ$5鮉8��4�!�4�&�@��Ј���@��y�	��$$+Hȫ@bg�ݾ��Du"@�`Z���;��Լ�U�-0@�8o�Գ@' ]�I��ة0<`����� ��
�v�#'y\-��l׶}!��0�ý�/d��R(��W� �	85���>؞���T����qqꄉB�+��6�㞤d��Σ�6A��;uG�4��B��&GN
*!xs���W�A�K�8�� �#����3�N�S�W�1�Pn���8�M�Є��2���S��:���Mi��4Iꔿ�,i�3��t�̵<�;��t�ǈ�t/G��m�k�vO̵�;���׾��&BU}�q@�CC3k���Q��Y�Ӏ�{B)P>�<^��������@�t�T��|'НC	f4a��]���ݙ�@E_CV��)�+�C���]3w�rkם!۽� y���M~@�kΑ9Q���j(�sw11�"T�$��۲cvf�u�	�4X˵��g�&����v
�.��;X.�NȄ~��T4pW��Nj'Pۦң�<�XZ�����3�/�2;�;�rŢ��<1v8�M"�͎������Q��K)]�2��M>���+��-��_�Y�g6�$߷.��]�nw��ҡ�a�ʊ�nZ�Ź�N;�=�bX
!=2j����.�k/V��k��>+�`!c��ҹ��O`o2�L���hby^�f#(]J'���7���t�e|-\�׮����!�q�m#�CH"�GF�	��C�J�)�Er��G�d����}�/�3��m
`�6��\����֏'�"~�/:J�o{?�Yj��09�42_$/w�Ff��e:��q��;X:�����j�ST�^�|:	���rE��+����W��:�z�'�.;���!�aB�t�聯 �}v
��=���[%�	}s������ �7�K(��5MV�����%6&�7Y��z��{d�}`(��xb�h�n�XJ�����o���_/����6���X����p�'w����w��1��×ٗPK   ��8Z�=�:��  � /   images/a3896090-6cd9-4aa0-adce-88a16a68907f.png��SLӯ�_� 	��	����;.�����!������������/��?LUW�\���S��"��A������ /���?���gl��@�� -����-=gΛ�)��Z�� D��!3A�F�kHv������� �s���1Cר���ސ��)�
��0�L�M �~��Sxx�-�[���0��1�:�4�Lr�<��'�K"@ $Iq ��\1A|�?jf��uѹ�#�� B���
��%����&��ڡ�x>@"�/��J#�@�_��>�ՒV��?3�����-�
"��>��D�v��/�_����B�����/�_���аW=�����,y�����K�ǫ�3���뮀�n�?ۜ>g�T�s���?u�jQF�dHO�aOüthO7b�b�HmE�����τS^-骚��u�i3c�/M��K��Y�(F-/`�Fݏ�	�7{_߽�a@��Xک������)��/�i�z	3���*�̉����(��u�{rq��YԷ��O3�D��Nɞ<�5��Y4�6��/�P>;�����N�컱oW��T0�v��g�����63��V����	��z��Z�JL��z��X����i�5Hp����y�G����z���`�w�����t��~Ԍ�zT��Y/��\?����J�8���3Kfd|<��Ԉq���:�r�=@�]�^	�Q�R��x�U���LB�g>�VQ6���?�:͚����0�t;aQ	���<�6��D��F�ſ�|'H�0��^s�|j�V#A��.���A�OoK���
��	������`��JL�-�)��1Q� j����4Hׅ�أ5͉�1H�m���-683_@P'ژ�s��F7Q�'j���a\6�ަ�9<�����O߭�8�%��z�{�Id?�ф������=]��EXg�K>�+g����H輦U��>H��;F.����c�U��{Y�t4Ä��A`�P���הզ��%{� �[F���9?�a�9ѻQ��*��s�YU$���̟.�x��9���ԓ���布��*����`�^v����tϷ���ߒ�p�ru��G@�'�V��dW I��O�t<:��Īȫ�Z����GӶ��횄�{�{�\M'ų�+Bh�TBTl Џ��k�%@&��e��v�m�g�������$[h�A7��>��>��~1=U|/���w���j��z ©�u�KX���W*
���2*4W�s�;�.�]o���څŬ����ۆ�w�)2z��>��/O��[��u�����5> �=|F���n��?���w>��R��	�֡�fWΥc+��t})1E8]�����*�Y}�f�(W�#2�'����=�w���Z���(��n K���YU�X!�&:���w���/5�e��	�r[Sv��h��΄ef�K�C�xS(?E�I8�x�D�SMҝ9�(��$m�h2�b� DH�L�A�fn�8�쩕�r_�.8&_i� (�?��ca�Ι�B�G���*�~߸c���a��D]$�j���a�N�0U�#��k!���%�|�Nw2I#'U�E�L����X������>�[����<�_�ހ�+l�޲�L�PP��ﲊ�Ez����,��]�ϒ��/�fP˟��C�vqy4�q�E?rT�V�:e���Eܗ5�C_.��ôh��pO^�hn<U+�)+��$�n�ט��0`*g���в~h&�ؤm��k����6Z��	ŃYh�QJ\,��؊�����#��������Oƙ��7mբ���޾��͝�m��.���Put�/����b�4{q�������@C�+1&�����T�b��^�%,��� ���2�돽�A�f$�J81���vs��_;/�B��)�e��qQ�<�מ]�l���F��M�23�g����#ޝVsz�I@�F�O�3X��	���o���'W��?��h�]� ����/%�6�W2	�����W��g4Ŧ�bɱT���G�(��Z4�jф���:�����Ϩ��2���X�8$.����5��GzhY	C���_�'����̻�ic�!��-���8ct�8[���Ʉ�j��%-�����{��hj�sav������+*ٶ <g�`6Tj\�O�Ɨ�^�_�����糪/��b>��J݌4Ht��-b���f,Eo�1�_<��O'1�cp�X�)Icp\��zF�� j���Z=q�9P��ؒ�V=�3&
à�d=�'i�]�^]5�+�It���^�)~8j���(@ek�� ��Q�и3̄�&[oV,d3-���Jy��%��b��J�˘�)|��DA��_D���3�!jNolvL�d!%I잫�պ���)z)�������/��W�|\���2}aH<�K,IY�Z:sX(=>���ZJ�HΣ`$��QJ_���BNl2��/��R�΄İ��򶏏[�fw�dR�g���s��&��?��Np���aS�����Fގ<1;��{!�f�c�8���P8��h��΋Y�΋,�I;����#�F�e�����݋%t���V��'9'@ǌо�M�����8���2pg�	�f�����˼�r�V?W(����r2�����5�(c�0�G>����BfN�m��J�0�Y�)ϫ͘�J�\�,AA�܄ʐ��1*𖌖�jܚK-p�����[�H�-�Іh��W
����?X:�����Q(��#�=�?��ܟ�����^�lr�r	N�6ER��	&���
����D?�m�K|�BfDw= ����6W���kk�l̶�;W��{<5�>q8h��A�lg=��Ƞ���!-Ni^�`{^�a.�^���써�eR�?x�&	���遘�}��$%Z��|��d8���/4�2b�����J!�k�iZt���ŕ�f����e��6��	 9����h@W��W-Trܣ��;���&}!k��� ��ݻ{�$�}TX#6v<�%������-&�Ĺh��Oo� xN��L���K�'ں�u�^w8Y��*;Ћ�����n�&���U���ݦ�z�����ݓ'?߫_��&�;��>-�x}�3��T��d�(5$�J2���ǁ�Ūŕ0`֎,�r,�����1�*
[���I����t����c{��3>�����b��|��M���&C�ʬ]k�i34��sPٟ��&ڪ��_j-�ץ�1�*>y�_�RɌ�ILD�d�#��f����4�0j�4勧BJ��!gF	��`���ڿ�4�-ؖ�% �ذ=n��W^A�#�}�6��X��\��4#�?i(���L�
�~t�.v��Al�[� X£_�����=��"� ��ݓ��4'U�L�Y�s�-�(ne���}k!��>�HU�gT΢u��p�{�g���#���Q�/��"�!����˪�y�лh�:�������:U���x0o��D��YO�.�y��";��El�ݤ�6��.�ߦOV��~ڞ��$��_�����4-?��W݇�e �a�kK�k�!�8用���==���t�ʶ���đǇ;Is�&z��D=��Oeq� �_�wrG����պ�U���Ⱦ���> �!�2�m�j<�T�麯����8ꪈ8��x\���vß+\;���6��^�2p�;v���R~��tGjs�1?"O��?i.+�$��/��
q����|ӳn{���ܘĿ�l	;��Y�d�B�6 �������$��<s���(Y�!�{�G$ (д����O��Q��d�|���)B���X�8��,����;�V�����یD<]~��DFGB�/�,J�O.�j)�gWWQu��^)
�4�sO����`�\�'�\�cZ?*���9֐������+�f����nGJ�㓲�4��Ƞ�,��֚[��8�>(sΎC�� ��|N��s�X��8ט4�ý�A��G����,(�x�y?\�	�-��~,Es��S�	7�S�{'j�#�8
�'�$D��D4]�	!�'(Ԧp��a@W{c����C�{H3�@{�׸���	��Xp9��k�Y�Й/��E��� N�A��ʪ}�&foZ�=�ȉCЕ�*� ���elsC��C%bXp
�\�Y����xr�"���6�93aq�F�7T����5��ci��i���M��!�\���Ge��Wf�w��rH��#Y�?*$���%��gV�>�f*@{Y�9���ra욅�kg�v.e0��(���cC+�χ��"M�9ܷDZU|�o�[��uw����M:`��@rM����;f�ٯ&%���i(͆�v�/�� ��n���bL?��������5�~�R�"d� s��ItX����D�6,�Pf�3�9	ʽ���i�\<��췖�=�lr]�(ڷ/�<�g[�/������4�r1�U6�n�%���͓��(4,x۴"T�i߾�l����b�h�l�hN�!��4�MKƶ��d�SNWO�x.���H�z�-p����+�\JұҺь�=}��!=Zcr�x�7����ے����"P�b�^<<�ӡ�mKw�f���Iѣ�Y��s^3�]���������S������������%��q�p�bg5l�C�n��~(�x�5膙����<h���ߎ�R��b�GQǡ�'rJ&A�r{rE�&|7��(0~"�G��V*B�S+�]]'ܸ���ZK-�	l&���wnhE���q:hҢ��ȶ�оXL��$��Y���D��ϡOQ�
 ��]�V�A�&Ɩ=�y�����w�ƒ���o�upy��N���[2��i
I���7kQ��Uf�tl�Ȓ�GS sP��:���ᆧ,G >�Bz����� ur�.˭o�m
���������U�V��jӽ0� ����G��<��|MV�񰣈��m+��=��A�G���&T��ʦ���R#�4??�����ǁ��M�wn���N=�Y$���6$X�js�C�c�ޠ�\��~�|�	58��+G������;
3��D�Q�36����h���vQ$�H�=cA�7l}��:�#���^���oШ�h�+��IǴ�,,���U^޸��<���H�au����P�]�m3!8S��V�#"����'��.�u�
ƫ'���TZn���q秪���D�dܻz6�P��t�BK�rHGzp$�tXjH/��I�W �	!�S�E����`�OG02e^M잯9C)h�%�K�1��í�����E���+����OW�MTV��<���h:h<�^�������}�h@����]�(��3�I
��?��+%ǵh+�O���>:=����|�
z?�1S#�W��>|��DR��,��	�9ol��	�x�I��ѝrG�TK�t�a���4���s,��p-ӣ�6�O�P.b���a{Ӯ�?�����⽟m��2��.(��~f���^&-�����H+�g�	_�N%��=�����>�l�u�|���s8s�U�._���@�A��踙ҏ
�֋n�nS�]q���1���I�D<A x�ß$=ς�����(Q��w�]6]CI��FHw�mu��F�Qf���]���Xƃh;��ˌ��B�4�>�(bRT&[�n����~��l߱?Nl%C��"-��%B��W��>�4����hC{?
���vNh���f|�1Ν��k9*:�GЉ�w>O�y���7Ѹ�1k��ﷅ��6�3�GKT����t�[;�7�9B�Ý�/Q���X�~���[6���m�3�FOEv'0j��=6?���b���]��C� �&5HYo��i�86��SB��|�Bl�^��Z_�)#��4���W�����:���w0?gە�<7+9ɒ:WC�)���J~dDW�!!��I�7���T�d����ic!�R����R@�.ɬ�2N��S�э�#���k<�H�ʝ�~9�f�
��Vi`5t)Wv	��&�-0�!m��:�)Z �z���-:��)*��LI�,-����[�5�Z�o��懑���N�8a�Y�啼6N�^�.?�AZo<~�	�T�>��S�����y+�'�z H��$�����2�A(�J!Zz�:)U�~�!����}�Њ�a��
�z�@IIyڊ�q�k���o��0�j|j��:w�旺+�V�mLM2�BJPu���q�a�݈kv�2}L[:�뾻�>%!��$D�#y,�̶N�@W�?���}���<�.9����m�-��C^�)2�u���4G~�Nxv�+��83{ ��F��D� Q݄��(�2�'X�I�+���6�w��D"P���{e�K� ��Pd����w�����t~��G�x@0M�x*��o��ܪ�� �x�T�����N��=�]�L:���wE�k�o���Î�&0�bl����{ V�z;4����=�
����F�q�������pon=�ۮ�l_f�+8R;��J/}��/��<����*�_7&ײc>��Y1%1
5�����j[�a����g�PKMߤ�`EOޛ�² fs��ZC)���D	2�b��T�Z������+���Ϝ�ǭ��FP�of6{7�dgpۏ��C�69<�1'k�r�#�A�'�1'O�*}k���+���ÙƾȦF�&V!�c�;k�o42������pH���������Ӳ��+���2��^cE֦:sT�}B���H��YW�3�I:##�P��0����yf�Hh�ŵ�uĆ��&�gz�W�H�Y���e�[��"�"��$�}OCi�<4:]�փO]Ĩ�	-��Ct�Ro+鞨F��޾K�R�gp�gPh��m��
�rK��� PU���GS����{'��6nw�C��w��@|��cE_狐�����BŪ�r:��R!�S��g���7<�q�F�:�z�y�yrL��k���4^}����v����V�$��B=�-}�FHpj%d�Z��o��k��̱P�fl#%ڕ���,�mZ��6��V6���W�H��<�!��_�>��5�;܅�T�AL�x�����.M$6�ӼK��b�]-WZڹN
/�&���p�*�h��Q��/6�sj�s�AlUK�|�C�E�+�)�Z4��Z�m@�[��N���F�๟3�O���ύ����'��
�3�1���y�gU�έe^�9����0E��,�㇉������U��Q3,�B�ږ�͔�!� ����" _���̒��hf���
��)V��K��Ѩ��/Y��!!������JL��pM����o�����[���v�ڿJ��'m��?	1�܀�� Q	��V�v���������S�&�&�dh�8�(����{ЮRpZU�7S�ɗn��^G�;��%%<��4�����;�GQ�C���:���7����"����-�^�#i5=�=�D�&�=&�0#�-�ԝAy�3��G�v1�`ƠﱑS?�B��=�ʗ�F��|/>E��r����c�Q'�k�+�'����xY�UC1z΋��z�e�\��6��%�i \����L���l��J���;*�n��1�/>vw�DA��>��3��}����x�����M�����ꟖŘ��FŇ4�~T�w���L���[8]��R�ͩǋp
V��d����b��Z�T6F���bnE�Θ��vi{1"��4,�������77czަ���:�(��w����%!G���vϕ��G4�\I6�Km( �l|��|Q@��*�[�B=�<�H��C?�_���s� �ɪ+����7����W��HW\�|��o&W7��Ksn7��<������I�h������s �h�儜a�G�
{,\�i��I}�0V��9{-[>��49�Td��*r�������r�S��fiW��h�IOܠk^�Ej�TV��E|B���v�z���	M��aQcꇞ](E�	Z�E)��Ê$�둞"�b��~u��7�9�=��e뚻=^�j`Tm>�n8)!wl���EyJј_�F��M��?ƍ� ��ZkM����I;���O�^�jN����b�?�����������Ȳ��e���t�nC��o����}��}b����S)��%%��V�l���
�c��+�m�������Ԣ��x�F3|��D�,�6.z��>ٟ���+0�[^�D^f��9�f���:|����Z.a��}�Bc*HN�X� ;QH˃�gsˀH��hĶ��$h'a��U#��S6��)���������{������>�ؤs�u�%��	�/By�_<���w]�� ��-�2�Rlf��ws<�]�@d>1����w냌��q>����j}H�S��2�Ѩ�d(�1�lBǽ�8�������Y��%W��h��4Y��E����~�����j�s�R!=�F.������Ľ�*�U����)+�J���K�rF ֺ�IOZC�Ĕ��М�!Wȃ���i�j�K�@y�� %�N)/�b-��`1��ϔ>D�Gv�Fy�U&S��$��=��Oǫ8@��5�(|�s7��/晗�xU���H�g�i�6��4�tS0_U������Tg!h��m�Nn�a]d�/�Ƽ��#�~d(�6��l�z�;�N��q�ܪ8�4B��+$���>�����ޛH'��~<��g�:[��z0:��\e��u,�9O�0nCUV8��s�<��~4N���/&��r߰ �+҉�}P�u��L�yu�ݹ�;�W򬚺&~�N��<��.�"C���J��|Vjw�W:�~<�H�i�#-�Xn�����d�|Ģ �V,�}<"6�o&V��r�(��[{����v\�f�_g�پ�v�M�$��/�n>�e	�JJ-�C'��n��KάW�s�@3����\��@޵R)��r/��f�5��HL��%$t�*l(F@��|0������ވ�"��g7�Oo6�Ҋ���M����o8���&%F��Z�Z)��,�N׎�����V��"*B�� ui�lO�=�D���l��s�/�
�#������8��h��V&z>��9>^�Τ�l&{X���adg(�a;�:m��.l��S�K���(+��aU�#曚�u��*���>u1,	�A��H:��BX_���[���J�xi5���TSI�Ս��3�ˋ�,���t�vV�F�	Ni��X����G�?a��i*`=�� v50�,k���g%TWr{1����:��خ�>��M �h[��?��1R��!��	�VVwa�Y7u��Ň2���g�I��8�_G��#<���G��I�[��<�>��5��O�?�\A��q���Tsm�6�t��(�˥A��ډv����ӗ=�
'P2���_��8֨�6]�vRˆ[Ex.���~�ݡAn�+��84�SN���r��ޏׁ\��S�۷@"W��X�sO������<� ���_���� �����}�K@z�0��2��D
��sɼ�������dA�^�g���퍕.�ܯ~�
����TB�3@����kc�^�g'.��^5翽$����z5|����1���a���F�:i�؈¸�P�� 1��y������ia�.@5���f���H$�| n�E�6<�%}��8̩E<�E�]F�V8 �vX��� ��,aK[�I�8̴�d�h��b�$�%Hʄ�#���GT:�A���F�٥��;?-��*�C�8yw�ЏEh��n���[�_9����]$ (o��m��ן���J��e�S�x/��esW?r��8�Kw����Z��uQ�z,�=�z��a2Y*���5L�P�/����%I����o�՗bU�o�C���B�a4�%�u%gR�wxF�uqK�}/��iWϮt�E�rTӆ����8���
y���1
"u����D3M6�@$e-�8i�.��>�f��bh�x����r� �9a�l�����q�X �v�w;pud�Y�2�ڞ�L�p?stn��7!lߥlm_GO����Ӯ���e�:���FP��(�iZ���Q���J������&���о��d��2��}4����Dʴ�����nyE�ny3��ͻr]6SUV�q���nײ��@���\B�q�Bn@쨒5F©G)���rU3E�}��I$��5A��Y�ۻ����	~��&kFǔ
M�	�u�J9�ꃡ�/�E�gE3׉��S�Ύ��r�����8 ��_��r=*�G�fqr�Y���A��J	�.예#)����o�Cή-ǯiY���
�x㟴=���`�v�1P��_\㜍��pc�@����u���Bݩ_h�4��C-�-f�٣���E�����/Ȕ�ם��{��s�)ݻˣۭ+��e��N�H���?g��O���:k�d��)
�H!�}v���_��"/�m��J�U���Ju��~�q[��]����D-e�1�G�X�́�a�P�­*ߺ5�p��{�e6L�������͍�WjX��i�E���U��������d��5z�ӫ�e���vũ�S+5�Ϲ&��EエW/���󈔘�f��1{'��ɓ�V��t��^,~���-���Y�g���t�R������"R��9ꆅ�u뀇X�޴m���R����S�bHB���c7:���_��{�q�:v��/���mc�����	6�ښ�ub�z�#r{.�{�M�`����_�?]�B�pN����n-���bGS�èv�b����BC��h9��-&ҍ�0j.�:�̨v#̼G:�:/��2������֍�#�(��35(1����x8{��/�F�e�� ��3��_�f"#a+]o�絸q��pm\��0�=e��[��.R̙)��u���%(�1Y,
�
Ο{�`G?*�1��i��S�q�����!D��7���P�;�X#5����ly46?m�"yǪC�r���ȸ�{|-`��b)A��A��¹$8�J�;���6b#�3��ݳmB�L`�5���cvNe�J���)�,�',MdP�˓j^#ai�}�Ŕ�
+ߚ�
��{u�e��T��-c�p�IPUc�
?�#�y��i:��DX�H�4�kz]r����Ylv�S����R����'WR���Z�Ĭ8��$�Z.5�V7Y���+	ިپp�=V�8?�ߦ����,7�-CU�.��@L��`}��Q��@���ղ�9}���o1�9�a�D��i�Ǎ���}i^d	���jZ��q�ÆR�m	�����ih�8�5�����2��Ғ59_�$�~'%l�D��6G��N*B�DZo?\U��j�y��P�yFl(c4Ŷ���A�|K��5A���Tf-���h4�YFl73SQEH��b��.����8���n���::�����#����8�v{1��O*eտ�-�,��4{����\�2=f(�n�-=��[��}�.�z]�coC*�²��gf��U<:0�Zt>�J�HSx������/�CUz>3�٤�K��������U��&(����ܳ�ran_e/Y��л�ee���i.����@
���ԼVg<[���_Cv�F��WC2��FsƏ ��֚di��fL
B����[]4���Řv�����v��3�p����=R��}��0�-�@���r�m%t-D�q�|};I�����Y��5׽�D��bS~��������0���\ߏd����Jiv[�$��O��.�_%u^�\Xȵ���v���o�k%���f�kj���ܞ��P��K[�"��7��k=gJܪs0�?�����}�RI�J$��m9Ƣ�c:y��>��6Qy8���0_1���k"6����-=,���'�����̵���D�����'�lqEzU��L�ȋ�hT��ut] 8V�P��0��c��!�I����pkf�K$N��6��VG�az*��Zg2�\Bey�nW�չ��C�GP���S�/f�}�.�����]��	V� h�T�R�je�2R�qϚ��zs}���V!3��_��!�(d:X��Z$�Y�!qC��$��a�+]�M��q�l'q:;�s�zm��0�Gf#WA�k�D\���w(TS����bY�c���=q����/wϺ����/�t��o?/Q�� �~��:a"��C����,0��t�`"���N�����xH��x'�},�4a����=�c�;p^�)�Z�jȁ���s�m��{��yi��������$�;�Z����};�$Zí��F/`��w/��	�]���;��"��;��0n|ؿ�
2=W6�;�6^	���v�@+�|�k����B~W?�ۚ��pW̑���~�r���]�}�v'���5��(����Y~A����,�'��S�~�ۉe>{�,?�As��)3dd�y�PQӣ��̯'�d5�sC>Yk��Gm�_��W�Q���l>�Ћ5y������Xq)�
5cR��z ̕��-qӑ)����Χc!���Z�q�jx�d4�Z�� �s��<r�����M#����8����0���+S��o�p��x��f�Ӿ*?����;�!�)Rw5�<����I��F����8�3�I更�ԍ�c�>���RD4{���Y<*Q���؆�ϣ��i�=�]�1��<e��wZ����N�ԫ͘M���r;���{�L���dG�����j�=`�T�����(��J�w���V��	�ج��b��Zݔ���RJk�so�|�	�R��l�Q�Ϣ���2��m>�c��,�Yi���Σ���4M��-Ǖ�2Ĺ�h�q;"��
�/��9k��^��7�R����� mR� 0�&�^�8��Nz,]��7 g�	*S��)s�P1��Y~�	��!��[�s�۽�30�$�wű)B[�7�Dc� �g�Q��C�:#g�GY���܄N8;�u�)�t�ہ:�E׵m�|�:5�'IN���@D@ �@�¹:��:�����n���o���zn T���:�s����c4�3����!3O0�%x�Y�Y�n_��>:>�l��������hZ�Q�y-�ah�
��t\v`���6ĵ� h�4%7�b�q�����\9�i_�X�I��kΩ�m��L�[����IX��0Bd���@����\n��<��J���[5{:��_�S�'�BH�@(���e�sSm�wē��%��@��q+���������a@dV����	�P* ���,v���0QOia�O".W+�j��,�R��+m8 N���8��G��xj&R��Z�܎B��S!,��"t����۝5�+/���+-�a��^���
'w	�[6�v��7��j,��L�r���h�2��S���ͽ�����W���ͦ��e���Y��)j>D ��&���c�/ �fm�2�%K��7�O������N��3�VF�>S����r�r���D����s튷3�p���1(�]6��6tQ{��H���7��w�"U"�U	)l}�T�ς��o�Ux Ch�eJ⠲{}q�X��)�Қ��ô>�֡o�u>�BX;{�ʏ�b�Ŷ�lGX3%�����!���DDs���!_t��Ɩ)�$Q��#�V��������b?��#��Lʥ�I�H�Y =���( �(�o����z���~�D�5�;��gB#��zDJa��(g�mϾ�	_�2�rC	z�㠕���/8�'��@M��\ĝ���*eu]�\ �M4씭$�լBz�M�[���0O8�;U�>���R���x�)�w<c��}@b��ot��y�÷4<fĞ�����g'�ˇ�'�b������4���D"�r*��	�W���1UU��},��AF��i%"oZ��)u�;+�����/'���h�	����L���~��Z�����Fn�� m8�~Ӊn�w�)"��\�-p)s���3W��}��/c,�#�@"�v�X�b �O� ��Y�X6Dɬ��1�4�!�C��:L�R8ct�ęrH:~L��/�!��A��+{fV���C�/�v
�0�v�P�G ��4a�2b2��]��cQ��dϘ�fqN�pQ�; �G�mJ�K�W8�z��l##w��O���h�m�޹L���v$]�
[i3˵[q�9�h) E:���q;���аj�`u0�ϑ�Q0c \�������B'�B��X��D�}��~�dK���1�3TO9���ίB]5��7y���j[�A�~mY���S�� �����`�&�}�rOL�ӄ�U��#o�~E����U�f<5["��wɼ��l�N��0x����r6�#�yϖTK�׈�wy�'k[� H����@�Y�Xط����<�6OG��,��wUK;`���,�H��O2�OC(�]�{����/��mSc�<�lǻi��g�ő��w�&?�ɔ6�G���z�/��9��@SqޥM,��~-4��T�tGPj>��/���!>R[d4t�'�0ΰV��-�<4��;�4���z\D�����0�ż��'a�]z�t>�-I���m�E$��\	�����#O�2��C��,�/m]ix:�?3��B�#ތ����|n
�bf��BWyw�I6?�kS�1�F���e�D��N��W��t"�ҝvz��H�D������ż&����$akCz�*:�UԵ�y����D|&]�ƾ�%�X0gi7g�cə����w2sk+a�_1�gϻ
���T[�����)��^iCcb�{<]�1~%���pݎ��`x����٢16��=�j�w(�j�����+O��S'�
��v��,ũ�h�36��O�����2߉�:����	{��Ya��	���WQ�u�$W��C�@Ўl?M(�_#@��QC�
������e%s��L}x�J�q&,�wC��3�"�$�A�=�c�w�{;�]<Fz�O���-T�G�L�o蓨y^������R�=@Q��d��"�	���n�������b��A����ͭ�^��?*����!ԕ��xzH�"�� O�e��E�*0\"H�Fr�ׅ�Xx𧤊-&:o֢��w)�u�� ؋��dYP[b����[��Fg�"w�o�卟Z���r��~���%g��6�t�tɝ6�����UE�|oPM�\쿠_�~F�NwFB�V�^����{�����;R�jaf)^��o��i�7�7���ZqΟ�(��~#a���('B]�����*�a�����C0ӽ�L
�{����F���_*H-޼i�V�_����	Y52�S��:�w_HMLg+a� |M�oal�<Ze�6�"ۈ���	b�"j|�(%g/�ź��qL��|�
4J�O�gMW��㑫��(w�pZV'Į�(�On�j��+S=�4�P8�oC:��v9�,�}rf����g�.f�"Q����Yφ�Z�`��⻔T
��.7ň?�ȍZv}�k�����[�����ut4�A��|��ڂɾg'y�4����O�$��j���}�B�������6溧�c >�ؙmǗ���{�3����
� �Hҍ�'a�=�MQ���r�O�������hw�!����������W��Y'��1����5��-���"/�1�H�T�AW_f����\~�b�;{{G/sJA��Ѳ�M��1m�o�;�r���"��a�ZiM	��P���V��_{��iRب�1ծ$]�{�HZ	?_��T�a��rj�g���>��_���;��ƓO�in�I����]h��S��>�,b 6�Q͌�����Rׄ�����wx љ2����/�5����x��)+2��1�Q�C_P�݅�J�#����z�2�����Bi�:щ`��b�n�b�)��pJ��8�Ok"F�=RT�G��+*	��,JK��ܤ�%��W�Q�4����߿�#2-�"�]�ǎ{Ʊ\��F��^黲U	RpU�J�I�6��E34<�8d��t���p��FN����CWS�v�}�LdDc����j�[1m��u�qɘ_7*�W�U� �t-f'[�a��!��t(]��z;�Hn7�β%���B�w��P�=��H��2���Xr��ޥ�'g@��a�fd�Ǐ��{����@a���+�N\�2��6�䆍aֶۘcp�͏n5ŏ>W�E�)�c�q�k����`�j6��=p���W}�}JF7��s�����w���h��dzJ}�Τ���?�&�	��8�+��VҒ����Ť�j���d=�]\:�!�SC�(��[�du'Bw������EN<�Vn�:��
�OZ�j?�*�*ח���koG�l�\I8���E�q8�f����q��>�������e�|�m�k�}^p�M�Ext=޹-� � O��B`�����6��*�y��j&�"i�T������u5�X��������'��:
�+��?T�eS���ܭ�)�����xqww�k�wk��Z�xpwww������~;{>�sfO;�F�P�^�J�ז3���i�Y#�L;@���Mj���<3��ŉe���(�wB��C�.7)�ٔvh��~��~ґN*���x���ǻ�&���F=�"=�J�ԩOW��c����ET��ǅ4�-�yJ�N�#zM��5��Q���U\�G�g��5�1f��5�J��H<^�&j[�-��`Nx�}�/��R]�g/iNg�/��QP�L+`����
h�|\,��V�R�Z���7��-��:��!�oL�qC���
A�Տ�P���$�耰'}Y�)�a�2�^�GLy��Ü�OC����ʞbI��_����{Yɤu?����왙�������j�q��S����\.8��S��L���eY cr�E�ߣ��޶c���A��� .p�c�4�b�o5��Ҍj��ǹ�=/D3:8�-����>7o��i�����>Ӈ>��qU�@u���b�*�W1(�'��xyX{���;V^�K'E���PX'��Oʹv��\�V�F��˪��
Iy9T>��g]e�◄Z,�3ޜ���d�y=��F���D�	
۽?){#/3諎�_�K�"��%If�ܦ*.���7i��}�S�S���b��>�z{�=W9I��k��[�e�m��:�wT_�
�+��-z�h��\_���;�|.���z��~�$W
L���ܷ��g�s�lEt�gD$E�S�S�u��j���g�0G�@�M\ļ��P�;8I���{�'4�^�D���(Bo;�x&Ǿ��T�C���>��cq��_Ll*��鐞Tw�2.�X���0��KK�ν�J�'����p��V)sW�<x����?*9� 8�z<���xz5x�%��&r��4�YM�4|����;1�����7kY>�����f9�nu�vP�d���یI��Cg �Y��/]�p�#t�H���_�Ƚ;CF���S���u���ċ!���a2u�=f@"M��ElQ�Ւ���qWNq�FyȠ�x�O,�Ґ�'��p��v,4yu�X��[�kOK/���j���>��U�u��� ��vȩ������%	���s�����/~i�m��$A=G@�+�M:8҇;��;��m��1ư.a�<��Zx�)EkU�({�ﴀ>�<m�B��qÖ���P�v/R�33�K%�q�*�M*1|�����&x�3�yA�5J��'�e*ӛJ��<�Q���.&�|u��,�������-�ū.1��| *4�I�bC�%4��߄D��>�ߎ�z�^s�=_rJ��x�x�0u ����r��ㅀ�q�5��ĝ�����i�}p��=42�XF=����������
=u\���W�h�-s�:r�m������$���[�R��[�E�2�����O���
���q�*Id�Ձ;MN� ӫ�m�2�n��ǔo���A|"�NF���Z�⾽8@��cT�C��}��PE�Y��5���^���V�r@�(�%��^���ι��	���j;�:R�7��A�$9���c��ө��D��I�e$�i��uڻ�/!�oZ�X��\�����U1���jS=�F^0w廋�r�
cE̽��z��Ia��R��J�S���/����a��gq������B$��.~{TXu�M�`��Ê�>��;�\�L�tܔ3�7��"�g��`���6�v�k�Ð�5s3|[%�%K���_-�7-��u�e�{�9V��ٻ��LY�J�S��N-���m�C�1���Uw7�@�C���O�e?j����d��6�9Is�&1--��P~%����C�G.���L'LsGO+����5ƻ3S�j-�����=#����ﻲ����n������q�u��n�'�{\��$|}p��ߵ-��Opo�a���Zk���@�����	��I�d�ĞN���8�9�D�n�	9(:�����@Ӈ���%'l��ȧ��&�;�c���@��1���H��H�7#j�{�H3o%͑`���G�)���%�ѡ���T�;Ow���[ƺxI��o��`�J3O��
2r�����#��G��,u�����LgU�����.�X�{~4�Kw�Ґ:��C�%��V�3�j�5q��&��c+�Ƿy�q��$m�!Z\%���1����+u||����`���=0!��L{��&�l �k��𽰼ߎ�����K]�DW����3���e�����S5�l&r������¾����m׻�]�b���~���{\�o���W���(-}k���3��_�ܰ@��� Y�A0���aB�C�ނ쏱 ^{��&������������?��-���bq�������p':���|w�Fq� �8d,_�*����(;�\�b�hN��s;E�o�
�HFD@*}�=��	=�I:ُ��Mc�F��g#�$��*OCp��C��@e]�u���D�T sN���=�?���z�����O�KC���1��6�w2�a������]�L�O���D4���g+4R�h!�/�]�+�{��ryRA��GA���M��$^~#�0Kߔ��HX�N�j�:�P]Yo��9�K�����!|>O�m��p��TxG�~���T`Z	|�y�,i�l�^r����m��6Q�ZRS�S����c[��΁�'��;1��P�sj��"�RIs�v�x���X�5�z6�Bx�������:)|�ʎ�����ydp2��x D��n\�B�ﶍ	~Ү���5 ���6k�ƫ�o�6�K��0��) {������=l��	a�Jg �)n���)��kL�4�
�~�y��d#Ny��Ѹ ���\�e6��k���xC����l^kQ��~h�ꮟ�p����i�w�yGL�L�7Zj���^��cg[Ň�6�(KK��&[���l���U��>�qz��[�,1�#k���b�9��7k���"��-q�Z�.��m5���I���p)m���pA/���$_ž�O�v�ɡ<�*�60� q�T��ؖMF?��Ft6_��P��I�����O9�yo/�G�m��������Z�����*,cSS��Ϛ</תޠci��Y���?+�q*��z�7���{@������z�*Ԧ�<Z%�*b�V�4���Bj�#tnu!��I��맣_���ķ���o
n�O�9�uh���r'6��<����t��h���4��7RI~e�%V�i�QE�����B��˵9����ɇ���Ţ���k�S�x��gV}��L�hTvXԭ˙���������	��҆�U���O����w���(���g���T�]t��3�c��vs�x�m�!<���o kk�y�C�+�#�R�Ab$n����u��	�ꄅ��'Le����"ߏ?��0:�|te�[��$�E� �Z��e�9(y)щ�����a���FX�� h�  ��e�<^��k��y�#�R7"���er�"<��i@�<�W��	{�-!mk<��I�w�g7]���� b?�(����[��r�Z5I�bHY:� ��Ð�7�>����O�w��L���z�����[1�t�]�ٞ�	8_g�K�d_��=JJ��bbF��4"6��(��5�X���p3	^_�	�+Sn,ؚQ�]�>]1+��0c�X&�����V�ݳ��k��;�dF�Nϫap�.�� ���t�5	<!N��A������=r�����M��mR��U��T�}����b�93����N�����A�N�����V��}6 ��Y�}�Z�IA<!�� �B�w�������B�w貄%�a3�o'+��;[��ϲ<D� x<���]>y�(�]��y-�"���M`��e���s�y���ήp�	B���?�W~�zޑGZ��}>�ke�tɼ��T]�}�[���!{͇�F^H�m��p�#/��m� �Ѻa�U�|�N N��W@��H��a�`��*���S�S��;�C!�6�H���WZZojFOLM��ר���[�Bc��]�to�nG���@H��E���ߵP,��1�.[��$�sQ�)��FT ���#�]��6]N]m1���� 1ČH�I���qUԻv��َ��ehV&}��,�2ו���ɻ,�U)�Բ�d�6��پ�AK�-#2���0�w����>��t99��:LYgI�i�\��ώ6�_����+��bn�妢��O3f.�VA���9�ˎK4v�
~�b\�2�U���^#n
�R�%��b+����)���M���xY,�iz���w?�C�â�x��
���fSřz��H2�����_Px��Ti�`��K�0蛜�C�*���ϑ�/������y���3>V�L��~�!�%CE���3'���뵰fEbPQ<^� k����}{���G��Fd@�o� RA�.�p�'��X@:�{
�f� ��
*�������fn�i�J�;ˎ�Z�$W�,	m%�la@D1��΂���&˒�uv�B�e�&ݳ�@���R	���Yҝ�'�?�ݜ�0�5�m�N�+�S���h�	�
$�Z����>�	����+ψυ�}�&9
��˕�~9{��!�M(�Jƫ�P8Z�;X��M0I�/@�O���A�"!FV��D�̍�3<�����)�B9�U2��}�6�|�~y]a��t	k
��j7E���+��x�ܰxtg?Gś�����������[�i9}۬<beeu�8��Ց8_W=��u���̐וW?D9��>fx�>k$�� ������G�"k�"1��K!�����F�����^ǩU���s,� 9��E�A&�Y�Y%�,�+���޹���܀m3�J�HqW�K�J9
�}
)GZ��Q�U7E�r��w]�[e�߇��i�'2V	?��Bм�֕���D���X9�+=��L��~˥sdU��8�s�ȥ�"�tԯ��-������P����n>u�����E�i'�h�k0N]���M��Ђ�\�����/GA&Xșe���>z�Ժ��k�Htß8=*K�� �����C�*f)������&�f1ϫJ�A�`� `���͵c/_u��c�T�eg�\��-�T�\�^���c��vT��d���W�7m��;9���g��"�D.�����03�1R�#��C��|�1-
��W~~�<���צ�h��v	����#G��{�*����t"Fⱳ�wB� ����!25�N�"(p9cYj��i�_ �Q?�c4o+z殥Ծ�.bK�|�����ѕU�,2U���/���� ��������ݥ�1�F��G��k�ΗF4C��p6h�s�I��M��XM���S��b�K����wқ�x�����8x���ћ������.$'S�B���M�k63�?(�z�6q��>ވ��V�)+st��N�c+V������L^��ŭ���_��)'lu��t�R=����!��|V��#Z���������͘����ۭڔ���f�m�$,ۺȰ�"ޭ�QI�jG��x��*,O�������7`�LyǊ�;���h��g�@�w���o2�������z��0=����L��Ug$܁�L��l�)���hT��Q¹����4����{_�� z�����H�#N��~u��m$��{����^8/� ��?%��asc���u���H�g��T�tx,��5�3��d���B/ySˣ�p>�d[�Q�*;+��
�fGC���ϸ�ZH�5?�/�/E���wqsyDyT��-k����z|�@���#��5����g���At���,�\{����d��B��_(q�M��e`�6��1C���qz�!e�c�C�I���������^��`Ox+�G�6gw/�pj������)Ö��̒������x���ʺֱz΀�F�+��i��b~���N[|�v"!�䋨�&w>�����/��z�PR��=����OZ���f8�]�D�2����"�ݎ����a������7W@�G�oȺ�+҉rR��N�D&��x����d
� ��v(󆫗[�j��B�v�z�[�<��*�ի1Ȝ�ԳR��x;�+z4�ݙi\ǁ�VJ-zԐ��MM��<\)�dda��*��~T%�_�Na�_�ό���T�i�x
w��/:wwN�g�9cp�hz��#16�'�o��hg�����7���9��2�����2RC����$����`1�c��pa�����P�.��6�$U+�@���r� �\hF�?�=�� �Uoh��E��2�8���@���W����TifY$V�؂�J���Z�6��-�8��,2�n��% .],����G#��t�@�5�"+��վ�`��{eÕvm�a��7�*G�	��~L����|�R�y�7��N���������T�Yp��;��ue=q�	�&P؇��-���{�R�4�J��5Zp5Wպ��tq�+��K�(Ə�L2

�bw���ڡ	�2����h�l�W�A+���i�X���&��Vp��Ã�/���ȼ=D��Z��Z�7�0�GjAkfMo5��OG�M�c���<��:r^��������tg��2��&�cץ�-#i�=谻�������sH���,�Ϛ���"�-͸�l�֜)M�,]��Yg"�[rS��g��t~O2 �����ũ��Zo3��Љ�C�a�c*�'���ܟ�+[��[]�r��#��|�,`ņ�(��ρ��eu�Ț���V3�Ҩ��>��<��K�����������ҍ�j|l���!�%�nGwdhL��M�ef<"ǑU*��=�� �O��3�0]i$!@��
����W�X"D���TQ8�jtCL����Th�F��!���A����^�����d��5Kh���I�x����J� ��#�r���O�Qnj�չ�:�t������L�ޟ����ʰ�.yu�4�b�V���C�c	�0	��I�W��'"��������Dn��>ڢ�˷a��q_Z���Ul_=�y��w�=���lg�k ����o���(yL���[E�W\�C!�cu����-Ю�u�w�r�g5��1��gmCn#��9��m�yW���g�����M�]����=�{��``�U�Z��-~�?$a�� 0��p������R{����LU��Yw����G��l^�����G$�݊�3�o�Y���ˉ���z���c00kd��ɾ����K4�U��r9�.]v��h�u�����Pyv
p��tAIz?��u��!q�P����8�K��h�ԇ����-�7��Q� $�ۦ���[�r�S��K�����Vr��4V���{�5�2�/Ɲ+�žhy;�]�m�Ņ��|�^B�o>�N�i�[^���T2��$Y-���a �y����O�s��x�X>�U��ĩ�_8�{�)�:K<+;�Z�JW(� gi���?�? %�֏{�$��F�~��2fx���Hh�a��5�K:E�&kn/�8Z{����D
c�H�x��`��
k��:H��L�rצE @鋏���H`%~K^$�J�J=]������@j��1��[��u��RΣ�uZ��k�F���Y5hd<:=@�R�d!˱�%��W��{�x�p�F�!���b��n�a�\t�~T��٣9�|­��;�%3�-9Z�t�`�����#�i����l
�������ի��[m���_L��L ��5�Rͫ/+��~�^�ЪH��
;^� ^���RV���+f�����l�׃�q�YD4$h� �F\�R��"�I'������&�L,�[w�Y��	����V���Y�J�p%��4�v}�0C�n1�H֛r|X�$w��u����-x#=�)�i�FK�� X��M��8�K��;��eâ6E�Ɨ9;�V��&uG�e?�21�����`�/K�@D.��2�!������|��XL"�H��	����F!�d�tB�TU����������-�W�QOh��x���'h� ��1����� �ӂ��|��Te�L�
7�ͨ���_�D:��v{�Ԝ�v!���w�d�e���]�0 ��J�u���Q�:%u�(�CƟ����D���]��B&.�_S=Ld}vK}���$mT�o���� \������2�`JK�]U�D�L��-�3����v�ϸ�I�#���1���wR���>&���zI��0�T����g��R����ֳͺq��^�˵���x\�IDֱ�n	 �7)O�	k�}Zҁ�0����)z�\9j��|�$%�&b^��~�B����M��@;�B�=ON�թ�N|�À���V<ᒿi�"��~~��i�+'����ť.�%�� B���}~ ��Ɂ�{�4�E��O��
9}"js9�δ���]5�H�k1��s9����
�����������m�@bf_OK�2-��A(1r<��T�����%�a��!�o�~`�����̯{$wP� +�z��{̛;��o�����N��dӅ�얫z�'}����ή��t�Γ�`�U�����P!'#�=
�H_�"�֩�,T�n�0�g8���̢_��x)��ͨ�֬a��N�De5+ȼ�SO1����f)���SŔ	q*��@���3�Lr�Ծ�C�O���yg19�pm��2���9�a,U��8�G~�޿��r] i��4�x��^۟	s�J��*���X>#S�|A0E��"ߦ�=d�u/iU=Gq�K�L!U��`.4��XQ���q�a�8����X/!�F|pˊ�@~՛J�K��w&��Q�]4d�m�*9gx�p���$���)#
ԥ��aʐi�Fܡ�!��݀<���(�6l�Q��2J߅�&ӓ����	J>\<�5��mEă�]n���U[�+�rP,��u%#�n�Y.S�����,�'�V�1p��d�D�鮣H�E�/�y�!5��]a�4�ڑ.Q�PFq~�,����QK\6�I�9Ԋh��gb���󤝔bxk�R�ꑰ�ǏM���LJ�/]�'�|�v�B{o~�(=rq�J{����	���yV`�O��j��!]��O$(�k���/���������c�l4�v~&P
#�4yX������]���)7L�eWY�͇�x����O�-HD�"�����Z�}����Q:�`l�keS������������8"$��8��[`�1v��g�&�y@��-�3yf��q�K����-����<���+���Tuݿ"Ԉ�cKf9,��iͶ�1e��-]�_�٧��0K��c"y㙄Y2�aAؐ��	���#F.�߼��y�5]��&>Y�	��/R9?ޖj72I*J�`���Je<���t��e�1��Q̊��к�x������|xuئ3(��_���Q���\ʊ3/�C�Do`�V4�o�u���F���ʷ�D[����*�dt�
!�dfv`Ҏ�I���X�����ޕ^ ��� �'nn[�����NF�t},�MZ]�%�-
��+����`#�r_+��.u�UJ�~g�J��IQ��d�ϣ�򌣎���[h��VH�=�-8E�-Y�.c)ڰ�0j��Zh-�L;�8��j�� w��F.d��8�Ss��q�d%A/�Pʏ���l�Z4
�(�*�c��i�AaI�I �==�[j�G6T���K�91Bb�^u*��n���4���+ְ����C�y��k���w��l������I��8���Y�^/����E$�x��D�HT�T�f<�졄������C_�S���t8r��H���T)�9����~���$���c�뜩��i�e>L"�Il�S�P�O߸#f[����_�����.�� ���a�������������<�,�jY��,2'�� j��I�;C(ڎKDf�-�B����ߨ�������'�:8��GkX��>���O1�����{ӱ�B��d�H3տK��_.�M�K���M\�O�G���ΐ�s�?ěo�QX՘W>.[��g�=�;��I��o}#5�O-F�2��	�KC�"��OA�a��g��&�赿Q����tM��e�o�&�ޘ/�ji�Z�c7�:��[L��	-���T\�ڛ�ѕ��m1:�����c�>2�\��r_K�^����[-�δ����Qy�M�|eYx�AF�ܳ���uY~�r���t5��_h;0�g��";Y	$�݅��x���	ky�ZM��	fG����؊y�b��x<>���I�����۔��I�/�L�H��yi�F�gQ�����-IV����+l�U������՚������>�k{?��������!i�����*O�8�p�&��fdUO<+uү���V�P���mݞ#����h����6ba��Yk��>�vV�sth,Ͻʍǫ�o��i��+M�GR�&I�v;b rȤ��*&���4�.䔇�I�^��P�+�{�g�C�bf�w���'W���m4���^I�ZŰ�����\I�"?��7����!m=����~8S�#���L��������f��w�������)`%z�O��ַ��\`�	��[V�i����D�7u�roKj�"�\�~�>'a�z	��&�^�n�-�g����1w ���Ь7{(Na3������klI��x�
QJL4��iA�Hw\[���M����)�u�x�ƕ�~��*�gެ�NM�08~L�˗h����l��!v?Uk�b�@�kL
�}��G[b sLe�l���3[���K�l����dB���5`?�S�L���7jC���k�Z�*���,S��.�G�:�Z�����-���!���Q̇#��_)^$���G�S�l�wi����q�e���	�'Y�P�����f�d6%ÖUR�)~Qe��
 �.U�&D0Ĕn����|/��g�aͤs�SCaaϬx��-�PY �!�aJD��p=��ט��a8�"��v�8]�vX�4L�1#O)��Ţέ#S�#���G)��h�a���g_�0�W��[�(êV�#P	����d�W��ے�m��o���Mg�k%��BK^�$j-5(f�6�m�~)���~����P�t^ip��u�=i�p���H���v�T��Z���T`ڨ[��6
}C]�B�PZ���ŷc��}ѭ����ջ�np�~?�d�Q݄��rd'�4�GT��	��O��*��k�c0�4�G� �-��E_*<���-������e���P9>�m�ef�&���ZY7��m�?����&Y&����͋�P1ľ�q|j 3H}�<e#b�7��v�|�~���I�������D��s�츴*\���P�ә�#In3f�H�]����c�zb���xz34��l�,��W�����K�lkB�q���o����~.1�Z�Pڳ�O��^c�+%mE�0�Sm����c$�>���c҇2Q�����<��T�S�bDR����a�6kd
��w�G����<�����b�W����)��,��˖T�����H����E�	}F-�!O���b&MƁY�������ɇ�Q���=���uO(MĎ���'���I�����$��V@.�����RB�6��s+ҕ6�袁�,R�@�p�4�(����Xo������C���{�]?�;̲�)��f{���h�:��L�c�W�3n�Ӫ���L�r������ժ�R�g����4�8�4J�+W_(���Ni>4f���l��~��f�^�9�a`�c�q�!��.f���(���Iƈ�5O9����~����DsU]�r]]Re����%=H>+� �#��+���3�;kN>(Ω/4�e��V9h�d8J)W��ǆ �F:����,v�LQA8%���@��Ȥ {�R�'a��ƿ����:�s/�Y�!�N�"�G�{� !���wM���Xu�۔ }$�λm��y�Xk���#n\�'ۖ�� ^��5�EY���d��������`�2����H��`�RHj��>�����4�pZΟá���nB_����ɋ���nM�h�DVf��|����[�_20�#u;4���]B�?��D|b��x��H�Bg'�s�ɤ�G* .3��M+dA='�g�d�-t�Smfgu{����_]bd�R�"dk`p[��Ɉ�y�Ë�ޘ���-�-�cU��@9��;��d���܎����Z���{�A�1������]��E[t���(���o[��{p�=B�L<�G�N�Eé%�
�����V�i+���;��nj���o�O�J���f��EC�[�&^��a۩��i�����=�,zi�,e��;ٸ�L6�B���rv�%Pv,�"�v��6[��ha0���?��E������Yļ�sY�vF\*��A@�����C�(_J]�"
�~�}�6Z����ފ鋼�:U��y�Ee�i������ ��s��s��sq��j��gM��"��_���otO�*2I=aU,<��őJv���5�oQߡ���L�1v�Zs�F4����%����\E*��phVF�:�K|�hɪ}{��1�mZ���t�3��a�Y`)�V��8�6��t]1[�Iچ���(���&��]��X���D2T̷�LK�c�ހ篭u��Y��W�-�і���5p`�G�9אַ��=gcv�S�_FI��sp6���ڤa~�A{�OԽQ8�!��H����h~f�F��[���P���kM�-�"�'$e#V:��{�6������8�� �}z��C��AB�[F/QJW���Uo�I�������r(����:�� 
z��u������ڿ6���������zU��۶'����``�h��t9�D�
q��e7htaȲ��կk0�X�(R1OA��b�����w�ˠ�6i^@%�ݰ���t*�D?5��/.%��~/�β�K�K���^��Y�]����ԯ� >S�ux/������ϔ��� 5һ�WD������߹����t��oIu�J�OYɣF����(͙~0�ھ�)��R%�VY������e��ЁQYZ�@��&�&v���$�5�]���jwv'L��e�t:��/�(յ5a���I����A�[�ߖ�ў>��gcQ�)A�
�rz�e7�*��L
_Pr�!��'Q�1U�{D�75��k���r�[���{��+��\7��$6.��E�/F�!��o����`����z����#�����$�
�ܧ���Ex#�,�����~'M3�~��6.CwЙr�+�W�gZ�ШK�_�����IlC�H].avq�(�63�]���r����h�/�n����9��`:�/`@gI:�^s�`R���w�����R-�@ktGk�3b����'d�Rc&'Y9v��@�<Zu���,�V�K����<�< J��<&%Hx�ɡ ���
%zS��j����dI��x�	 #5yN��7Y�m/(wx)㫿�0��Dr.�≚&�@�`�)b���֓�m����x=�
tX[D��F��^0�^o%��xi��������?���`8Q1���25t)R��D�<���4�js���#p&{���e�j2�0u����(w�wɊ�����Zl*��}M�>kN0M��U��/��'�|��b��2eM�>Yjbo=�_D�f�d��Oe �BF�tBF�@r�t|��#�7��M
o�)7����r��p���-^!�����Pϊ4�ѿgM	�)����1�����0�μ@����;�p�����e��n`�|��.�(v�@������P?���>BRZ�L ��m2�fK�w}���m [!���UPZ$�ү0(vk���_�IK��X^�m�T�����eW��ד"�R����$|�Q��U�4XW�� �{T9n�Dao[�����ӂ�)<􎬅��Cj��|д����AE�ʏ���i��U�<�TPt��/s�]~b�ci�r&�6Cz����F�݋�M��N��p��lw�)�T7�n�*��q�+:-l���U��+�J񌴫����K�JCI?�~)���%�|v�H5m�����>�Ŝ��cTm��8fo�{|?��nziIg��D��2%��N�@&��Xƞ�iN�mAu���6�z���{�~�X{�w�x�x�X��:��:kF�; �q��X#H�{��#�T±F�)z:d�*�9��52Z�.1�?�5f�U�_f�ʑp�ެɑ\(Y>M��&ǜ��qJ-�XV������zJj�/�q��O�l^���Z�H�2�����^B3��M9:�p�,-�v����2���*����e̝���Ȟa��b|u��#�)ճ�S!����}� t�V�����x�@MTS��	�R2=��]�]ί��Q0#˟��A$L���7�e{s>@zVó����q&ex
~���)K���5
���Z�o�&�u���x2)Ocٯ��pI���e��1��~�7�?���!�)%Jz���ߺ��X��%��3�B�vp�e߯�'�P�TZ�|�YO/�(65KT���0?y`�q�O*	uj����|��mN_�|+��s���N��O�2R�B��S��;~���̷<��r߶5h�!����x ྆yc
�����:��5^�W������v��}�{�e�����b�ˍ����ƌ�=ai���S+.. ��]�xnI:+J\����� ���r�3���UA�V9��o��@&&�\��<�o9���&M�惮��}���w�d4�۟����ŞN��l�p]Ξ�`�@XOղ.�φJ���"K�ǍJ���>cJ��N�K��Y�ә������|c4A>?�N��׍��ա����ڕ3�Q����N��D
s��ct�g�k�7��r�L�f�N����haV�~�^�������y�[O�|iT�
6
����I
�}f�P_���K�F�W;w�Jc�O���X�_3Zul3��ԗ����*�u��a&y��w�г�Tf�z!���4���� ��x�ۨ{�3k�n.�f4;D���z÷�O�c>y2YH����Aݡ��0�694Ʉ�;�^�s�ǭ^~�]��vc�H1�
����C�[��a�|�J�L�=��9X:q盽VW�V�Ϥ���-3���B>\Cm�?x<���Ηg�<;D�1��|��qvN�H���8�u@l?1�l{h�60��#��򍍥���v�3\攳mTs�'#T�a���<���n��^�����k��{u�&v�J�wvR�/�}����g}�����_!:9��n�D<7�>���!���@xx��j�[X�������i�� oԸ��:��h�a��o��e��y���ei�+�:�����i� �f����<�>i)�k 	SK���[O�-�e�6��Q����C7��+�C�k��جZfNH*e�2���Å�؏�k���	�
1�
/P2��\z�{2�3Ӽ��7�Wc>W��"�����94�=�4����AK�,4����I���&�lV�C~�[$2��평(�$K�֣m����V\���2M���b}�џ�g�J��v����+\ٚ�H��88��T��ʚ�����'m>��$�H~Y[6�Z�Hވi�Wh�(���º�w��4�2�2#96XC�>���R?C���G�4T�I�df��_�$�'��P�nQ{�aT��<�%��|�?�aq�����ױ�$� ��ߛ{KG��o���'M�?�r���/9[�,M���g�+���sK�����><�Y��i��p٦"ݢ�&D�{S�QZ�Ն�LsM�ް/+	i���R6���dk�G��.<?\���[��ſ��:/zb��0w�}.F��4.f��ӆ�dq�YĎ�)O���C�L�HF��TE�zLb�)-Y@�s�m��FPv��ɡ[7/8�w�x���s��d"6�"�y�2�?��"�<�BW}���2�K;m��Pg����.CA��<O�A��j�bx���i�/���f��i�2��TB�J{�gjt=��`s7g�e�-�_ ��i���a,/��	����;McZQi����"]e��"�������o�8�v �-��h���Ň>ēK-`f\����$8i�u�zsU/��T��cS�%��m8��O��,����]�x�R	���B�
��zJ�yv���uF�����'�YA��mSA��v%��q��3�)�X��\|���J� w�������:���J\Z3T�m��_�gt�2�Ϫ�+9A�G��ɚF�_�U���()�Us�^��-��
�%w�+��ޒ�?.΂)h��� ��Bp��'���6��!H�������{p\���S���?aKu��{u?Y�Zuj�땬Tv�+;��G��~��3�2H�U��=�=���"`?G����8r̰[-��'�	�_��>��q��=b�� ��0H�&>���*8�S�籤G:��:��t�+�癔�O�:�퉂��x=�3�s�Z��K	cM;o��������K/_�$9+�r3���6.֑Dkֶឫ��a�:|{Ī��贜�^j_��8�5��ѯb����R���.�a���8Wc# C�,f��E�~����߮x�.xl˒ܱ�D.B*�^ݤ|��$���o�g��Z!���� Q�y���
�u�
X��y{C����XF��B�k�R�)W��g�>*�$V�!Ӑ�+���"5)ٰi�\�bG���`z���|�����׵��l��r��x���6�Z)��W`F5����D>[d�:w2��Y,�<G��,1�<��(����݌���>������KjU!b�X�SL6�P�~2R�/H�É,Uo��۴�b�'�녞�i���Luxidf'ld�U���()�=L��4PI	7���6\Y���:��ױƛ)�c����[�����������\��9w�|"k�9`l�K�:Ο��k��O^�!yo�-A�O��������O��r+$B�M�8HY��>��,]��3�#A���]�5z)Hu1��Hz5���b�Pͩ6�6_�_����oyۄ�W��=m���S�_�h!��z�lQ�^ !*�v��g������Wt�%�[�Z���q�p<|�ت�8�M4�s�T$R�u\j`˃�\m���>w�8��Ϡ���t�6Eg���̠ݬG?||NdW�j�D���RJ��vG��M����u�����X9�������=9������9��ǫb[�(�437���(����n�Ǎ �&�oG
s���5���Y�Gi!�\�PC�P1���!���9X���kS�\�V���^p�x^�O�Ზ*�A��O���f݂�4��L���ʾ�el��mv?�<������l�Ԝ����Ƙ�ѵ�(���gH�_~D[ʿ��&n0������ݱ^��c�G�@c��»�Ёm!f������]���>{��K�G!v�����BuM�X���W��-���m�*��Ʈ/f
�O/>�n��,Rc[�'���7������w`�;U�[�a��=ͻ���Y�a�/^��g �Y�V+�b[�r�2F��rxO'c�J EH�����@*F�8��.�`QX`�\�XLG ���8Bz�Go�}�,OU�1���DP�BnA��I�`d�Q�����MvGD��z\� �r4����K�nPQ�������C����y�q�>;P�H���P���ϑU�XE�7~�f�lTp��EH�^�mh�+а_��Y I4����s>�N7�c���%/P����7�$E-1��1�w��`���H�p�<sιW2d��X����8_��p:ڸl�n��%�&���w�
Z�~�Z��H�!�ц�b�k1�՞ܕN3�����,�	>����5��
x-TM��?�		�([U��U~��һ�VabYG�Ref301������u�I�ۃ����������Ϋm;�R��/ת�d�н"�����煱���;6��k�8��3*�9�fr��k��j�X������i�qL1$\+SY��D����"�Ū([e�̂~��F�ft���0�o_����Yn_F��1�Dɓ<��߇be5����F�����Qm��	XRV�����w98�-@��2�]'zйwŢ��M��1�27��~8�5���`�˸�|�s��n����c�q?���gu]�O����2.�d��9D�������E��l�b
�}cνӵ�;�����i�G�ӱ�ɚsOw|��D��Բfk�c���ch?���tB�9v���� g�S 2��*6#�	Ë�+�|����UC�?�McS3_c��7`xi�8�i�zP/hw���d�F tr~*�WE�7�PdWY-t��h�߇c 7U�_D�����p8�A�1�p\���7�[�3�ԅ}y̥�"�v,��Y��M�������҅�Ǖ�@��293Jr��Qa�����L
��-kNɘg����1�uf>�+�� �J��s�@�0��q��t�a�oo����h���T��to����1�r9W��>�9���w��iH��4[yӦ�c&l��
�oP��AfC_YD�
�h�KKىq�#�d������i)o���]ͱl����:�+��sp%��1lׄu����˅��s҄j�V\��_͙3�:z����!ԟg]o�f��%`RV�&�U�m]�ʌG�R���5ñ��%�T�[��������Q�I�B����>����O*�W�(��Z���7Y�׎xb\&��Q�L��S��5������8���w�੨�ݽg������=��aq�nh�U~NXU�C��)�����q�n���a~D������nr���t� �y4��wi���A�(��z��I�ɖ�6��QQvv�	��J,�������:W:���0�q06�_+��{�@B�<�K	�FFp�~�F�〫��f����_��l�?!2�@�]lۣ�[�hT ��`X$�w�c2��/�E>r����̳���@9��e�Fد�O�t�y������mش�*	E���`x��j����	����e4y{}�Q ��fkt���ᙬ��?�-|�C�p�ޡ��r��.Sz&bBA��1w�S�,���}��B͋fx�ٴ�>��i>�G�M�7�_�J�(7`�P��,�I��EO�[Tkt��y�~d��F^�����^חb��˚�DS�����iw2�a�c�<��Y��� ����r��U�_Bސ����y�����F-]�������a}�䂙`q<�%��TN;���L�#�A*/�c�J^]W��@�?�d `�O��Ƶ�˶^:m$�Λ0?�^B�/�i���gu"v�2!���@u6ms
��Y���2nK�P�ά���e�?+�N߄��ٕ����}P	�1L������� ��KЦ�4tQٙ�����~���`��~�og�5i�ҩ��8R5+��XF��caـZ[i��QŦh׀��Z��l;��U�(�2\��？E,4@�oZ����v�O��̎��vElIw�K9�Lk�o`�H�w0�ϟ?�̙�'�'�k0~}�����`H�mM�f7���5�1�{�eq8�������}38%�(�r�/	|r�b���2�Wu��?)��}8�@�[��Lq�e�9 2�*��s���r�#粈i� �I�)��$>=�ׄ��Y�}�߅�u.ĵ�\ƷL2���κo�I�|O	-,����L�e���1S��05lt�́�=1r���߀�PkM�l$Z��F�E5#�	ܚ�̊0b�$���G����^��!ZzÔWX�&�!�G]�N�c{$�����{-p��U���}ڱ��xz
�ݗE�x:<��r��Ǻ�wF����a���o;�2��{c�g���k��v�q�ū$�@1�"�\��=ɛ,�Ѯ��A��>~�Ρ߆����8�͂E����i��̱uf������>GX�gi����eh�)����ـ�mo|��-eB- ��h����'J��s�Y��?jvl�e V�Y�2ix��&,�[��5L����PG�@P���{wk�w=�PK�F�6z)8Ԍ�n��N��x��>�}i""�i��;�A���c�� m����Vh��C������&��h������:Y%����
�VU�Q1aZ�ϩV\�#�����8�Z��ߤ��o�q�q~C9�lba�P\&k�$gk�W,Zwߐ<2Ϥ�q!_��>��ݰ%�H����6jL�f(�^O���N:���p|�h����˚C���І���p����C��xPJ���Y'�2�	�h�X�f�D��L��6m�<�%�P��%Tt�-%xZ �h�db���l�-�':������d��Yx�ZW�w��AlxH����p�����)k�4v�j����eK#-1_�z&v5��� �����u]�ˮSyCŧ1~%^>�W���ױ_���װ�;z�0e�Ĵ�O�g�ݯG(����߭r�E�?�oa�oda)��f*�ֱ�E�nU���Dَ�M	S3ו%?��]�b�%?L+���G���QQ������z�<_����wz�Z�7�Q�І�n��ܡ�1W� @���9�����L
�45���������� i�ⵙ�$f%-�`r[E�̚mɜ�;���3��c��	����͹(Ʀ�S�1�k��f���+'o�':=w���R� �Q�~o����5NR*�
T�3&͢+������2Ź��F�gm
Y�tn}8Nә�ّ���<�C��ɢJTl�_Dz[$�:��]�H���:τ�V$��w��g�ܳ���Jyؽ}���:����锥���i�Y@����B�L��g(����C	�&�WiY���u�#�i���s��K^@CCܾr���A��~��R�QdP�j��;����aƳ�r:�Qe�|��%&c����ǈ|��s�5z5����y"���wr�_F�SD]k�j��ũ�e�|��輐3�X! �7%�>���aK�గ�-9q��_���J�>�h��<a��d�m��/v,���Ili����l~��3͗Y3g�U~K��{~��`�On��Ͽ�.��}+���5�u�NL��_��"N{\���ڄ���p��5�?����duUАťMY �f;jN�L܋&�V��M*tW�_ee��wmF��s�a�c�a(�i���S�E=��U"UHڑ���euT3@�>ֻ:MuԆ6B'��k���W���
�k�� ��~h��
�[���&}9�����V!0�+R� 5��"#��$��@�nT�Œ����
�'���z=P�I}P��d�Ҁ+�ȍ.�Fq��V�a�}28|�P�a���SoL�u)�S�P\"e�Ղ��tJ��)'�B<�)�����[6�� �H��kv0�/f�ll̍�xN�x1䱣*-5�"ڐ!���uaZ�;ks���>�~106>1*�V�e^D�5�~�Ȩ�ԋ�^�����(�ŀ�=耘�B��`}-6�FX�k:���:E�Fdw\WDNLP6��	��8��^ @'�灐�<��������4S61 u�����m����+f�,X1b*U��H���] ��U�5����3���WTh���Pn���a ��R��A@���m�=m����8��g�|W�rg�UFS���0J�MeB�D��nq��J���ic�I��|�
Y6��~��{�*Vα�U1�����\a�4?��CH�C۾���-̯���g|��M�36�ݾ[WXW����'X�\o�
��7d�dJ�����a�ҧO�g)��VV'��F�'<Z�Á��&�e�� ჿm�7��r�\��-vs��¸���r.}�2Q�t~e�%���D�1�����D�xc�$o�@#ұA��6��i�0|�E��a�4k���I#�N����f"��%����W���I(�O3�r8��� [���u�@��'�J!�,+� u��p(n����>/y��-rau�oȊLc��Qb������K�<\���MWsU�a"Ȑ���t� �b[�|0]~ɔP��88Z3T�S���vY�\	X��ZUkOݠ���.؎����\�4*G�P#��Lq��V�+��*��������ȇ�v��U�� g�I��'_G��2&Dm�bVp�&�A$��j��e�m�2}ʋT(r��7	1J�ܺ~qm~J��&��	^�:6�;׷:�LR�b27��P]� OX��s�ށ�&��X�Eg4K;m�򿘜~����>D�A���W���$�vmW:+.�>h��P]	�~MO��1�~ݕ�0�q���\ҽ������"(���ߍ�L'��|�=�;�XG�P�&��%��X��,�����n�d��wq�|9[x7p�]��~���n�+�q��n��ñ���S�-�ׇ�T�?��jk�q]�%L��[m�d�vV�ҜzK�b&N��ţ�TZ���\��ѢЮ!�C�Mа��$g��~��N�\�^�H#�ܟ����O�$�NDR��+�i�O?�q%Q�����W����T1���ɚF��>��"O�u� 7���~�=��?n٭ƈ�� ����,��;@����� ��:F�y�O����z��j���	 a�*��F|�j���-o�G���n�a�R��fr�XJ�J��o$�����Ө�<���>6^0,�*xP��g�#��P�D��,h�!N�ۦG�6|r��?�a4%?�/�<N��,>{�댞`�#��0�A���o�Y�l�j1���"��������Cĉee@����:*@`�{X����b�*�B��U�b�q��V�Ԡ�'ǣ�>�ҙh2сV}�a�8I��v$�S��GH��4G#�j�mQ5�j���*쥲�w�ܖ�����E����=��ousI�A
Y4��hq�n�en��?n�K(�_@��u��-����h���C�խ��4zXj�:J�����g5����p���w��XL���������i�񲢗��7�`���7i�ykd2@N�Cs��@���zpm f@�6��Z�%�s��	7�Su5��ylND��{y��ܴ�Z���*C�=a�h 2���f��X�z��:�N�"��t��ͭ�F�-ݶe�T��af��Q����R�a=�! l��y�����/���&�ӱ��ޯ�+=�TON`NgxW8hV~�|��ˁ���nb��3^��?�P�uW��!����Ձ�1($6�\�Wc�9���~K��32T<�ju��Τ(w���L��-v��@��ދS� @!5)JA�V)kV�鼼�+���kʧy����(����W(����a� l��S'��뷛��M�SMC�����!�͆��� כeh��ֆ�I񏳗�7��M�۔�:w{��-��T�^>hm'���>飛��S��I��sߥ$ ��:u�:7�1��	O�$�[H�-��L&r�GM<
T�R�,V����ڠ�bZBd�������RI��(m����]�����<!} ����v�H6f)����L�"���m��5����|��E�S+����hD�����M Z]f8�>1�̹�i96M�x�bc�!�c:�L�����0η:���|����}�� ���_6&k(��.fp;�R�r.%@��C`��n���L��x#mV�E�[����Rj�;�h��� ����>/E��E9F�.rK�nӃۺ'����A�B���dl� ��������p�>o1�%��"Ęy�o�n!*L����I�Z�> W�[C�SȰ���"g)<6�N��������B�w�y�i4\��3�Hʹv���Ԏe��ݟ�  `�ngD�@ k��EtC���DI鷋<�2�B��jd���g�r�y���[QݝD�/=�?��}x޷�^��s�W#��wKWS-sa�C�bOG/|�O�YD��5c��_Vo�K_^T���5̗Ĭk��@�P$F�}M�N$�<�By
K��2�ȓ�J�`��R������
�l�<��L_Ύ.�6"����.��4t�yݔlw��|Y~���Rдy���|`"����0�|Dr���?�2K�,)8j���5�$�vC�z<��`m��Bt�[���p������S��B��Ѣ	Cs��m�4/6U	���T �ET�2�V.#Խ���ʳ����u��O?�Z)L�^<�D�r���z����~
��� �vܾfV��c�':�]8�Q��O!���w!��Ԡ�h,�e�We����s/~;[�m`�0C�96Q�,��6a�7f��-q��UX��{��ؾy���(����5�Vf���gN+��O��]e�#��4�c���E���)	`���񇸪%~s���"�c:KZ�c����/H�;���2�uF��?��OXl�H'Js#��й"� 3�ry-�P������NI��<%��m��Me�����cKT�Ap�ݶ����+v�����PF����m��]m1~�����`�b�f�<Τ'f7���jӼ@7u(��鎢�5�h�ݧ�������0��mŉ�9����ή���^�k6�' ��g�u�F�F��;z�����C���̧��sZ���y��n?k�Q#���:�h)�:���2�"m��YL��oI��GW�J%��&�����zt��I����n	�rE����\&~ ���DQ{QZbOh>n� ����#PWb��Y����:Tѱl9�o��8M�[>�����"J�y��Յ�T�Dfn*��N������mZ@�d#Ď���*T���b��Mo�b����V�6=��l�X,�C*����N>���`�U��7���S��������,x�ԙ�(M9V׉�=a�!#�֜Q�P���e��g�bs	D�[��R������^���0�m=�=����]bJ�\��7�B7L�;ΤH��${ �x��`�~�!��<�ۺ�d%�'�a{dZ��@[ɆoiɪUֻښ���EGMa��	���["Ѱ���P<!�����F�x�?r�䭦�AR#�����%�4��)/�ʠl�0vY�bm	qLI��~��odW��{۸Mkw����?��p;!������b�Ф�.�v2oP���t��>���(dT��A1�?����8|#Fy�Ќ�U�Β���gW'�|W����/o����l;[��t��c|��O�C5m�2���+�A%BfǶ�y�J������#<I�J�sR
�Q�,���q�yk�W��r^?`P��߇�{���޻�����Q��mo����%�v��J.�wT�_}WJ�(���5wڠf�.�} �P>�J�r���*�L'���G��ɯĥ�m-��)�s{�:�����G��H�9��4�}��}��(l�\��%�D�5�%�l��\A\-2��g ���-q�[����@��;��R	'"��Z `SYQ�{:�{���x�ȥ�I5�����oPk�>��u�w&iΖrn5���r�965����aW"n��:j���J��φ$�)&��ʥ�N?!�Mkx8�[ w�̞��1����e��EL�.��A�G{Ӷ���r���S��*���E˦4c')?���KS���D^~�����t�Y���;Ȇt/���o�U�mx�r��G�Ĥm��-��U�G�����/���CNC5\�c����O���P���A��S�ک��q�T�u/����6�"�ꜘ��4�ȏ���7|�^:��g[[��j�x�ۚ����^l�^S��G��wЦ�������7�)��U���l�?�s�]	Yu1�k&(=o��=��V����:�%���ˮ=�BO힗p�p���-���c��b� � 2�ɮ�s��9�*n�3>���}�&�A)m�B��l���r7ESA3�Z����]��d[ɯ��m������ܟ-�q������0P�%,7��y��5F>?������6��%���B ��;���
j�30����ߦ��\��/s�����o�=���6@�yl��\���}pq���ƕ[PmX�2 ��P�. ?����i�o$Т`�I�qD܌��6��(�����Ȏ>�?����$�K+]9@�Z�߃R:ڰ�F�+So�A�ÌB�J�� V�8"����,��ϑ�K-^�+~3����R���M/����Ur�;C�ר��Q��Wĝ�'>�Ƨ����(I0�m� A&��25X��w���l_�cVC�zJ2���i�M<��w滙�JV-*����Mgp�	�0��W�4�S����v�u����F����ǿ;Ij�_̈�H��*�v���*�T2������,����c�`r�A'ASg3�\N4�H�݄�t��}�\j���_ջH��ew�1�}�U�Fj��L���_��힓�ޖ=�$J+ded��^y������\�Ƭi�+*�^�D�V٨%ύủ8�\Q��S�6?D&��=�Y)-�C�jx��#9��˙R6ȑ:&�Ʈ��p
�kDj�9|V��+ј�t�
�wfBY���JQ�y�e���t�'b�[�*��6�@v�J�Pv>�@(�|U���� �?���h��A���z=5�2�Q���� 9I�N��yZ�}�M���>��v�i}ʐ��uWȺ�����~"�Bj���W�������q�}�Y�����O	;A-�r�)|O҄tՕ�eQ�����������~"��q$����U��1���Y=���%�GĨ�9*М����(�����VHc��l�u����e��α_�1?�� �/f�`5�Bmd�c�_��b��k8o�wG�.�M�!�N�B�`�6!�P6�H��ֹP�wi&vN�2HZR��
�6�q��L��lk�&h��KI9w	��9O�?v�z?����Ԣp��Ӽ����>k����I�{���Gc=�8��ׂ-��lcee���G��)Wa�zן����Oɦ���I�e�Eq�J���V��d,�T;��VnBD.'x����ͥ�ҽ���P�j+���5_��'��s	�O�lB�y�A[�=Yc���>�o!z �3�x/�^�m֥����6P��9��LС.��i���A��]F{�G��H@����p�.��蕾�~��RK� Wzq���D�B4�휳5�i�*M�m �R�lH�o���(H�%H�2(��#)>�	��i��"��t�x�dk/\��� ��׺�V�cwyi�5Z	-`N�a=����ѭm��F��GYz�_Ʌ�"�+"+��3�bmJb�"9q�M���t�h��麟���<1�!�l�Y	���_��3��b�~l�]������65T��T��RȫQ�����{�$�Hｾ�銄��)?�T907���fq�o��⥋s���v22�k�)ba4[
�QΝ�a1�#c���>S�,�;�B�v'�3#�Kg���3�tCY(����U�d�X&���gK�T�
wS��_�t�Zβ�P�3���,�l0E���G���!S�j�Ϊ�3�V
�z���[L�/}ﲨ��of�Z|1�}\l��~�� �Ot�0���Wh�J=�mj7��v����%�Y�R`�h�-%�ӮknFdxr|�ByL�XG�l�����X���|%Q�=<�O�����0�xmT%␃�Xv`����Y��c�B�*4�-'����o�젼^L�;��y���ն=6�oE�0{B?�{���\v���ݵ�Y���4'�k��}���Z$*�9v�,�[ʃouph��b˾7��E����w]f|�4����\��X����p��k��s������mX� �#�E�S�f)�ϔ[b�Q�9����M�S>V"M�d��T�>���F ��B��c�ת�x�W4*����c����/Smp�h`a������\T���ᬠ���/���f]-���i$=�lP�̽V��Y��T8�~��u�ܧ��X/Q���|M#��>&L�%�����p��凐�=��lL`�צ�0l��#�%فe��b��%B��\OW���1��0!�t�M%6�(���E�dTL��/Y��)���3Z~,�S@�KYͽ�u���N3��& iAd�[���b}��00�X��)$�C(2��/2lE�*�F�,,��e�����n��K�nr����PX�O�+$z���'yt��K�h?�x+I�7�P�6�s�)��J�NSG	���*/K�i���%U��0�n[y�WS n��Z�� V�rM\6�1=}!X��>��ʨ��!c�3Pj�ف���J�;�0U�=��S�ʺ���bw^q'B��c��pf���f~��i���w$Qy {,�&¦%j���O�����G�ʑN>7��NOf�@0��H��'=�%�8���ѩ�$��8���]2���c�Q-T�M���y�|Y��GM������tf��� ��(���[��5pH�$�:Ya���I�#�h�9`��wl�U�m�L��S?��vo�GB���*�f�0-�8�� -�kJ.B����B#P�������!е:��r�im_֬�F�Q��1��=����0�R[L�xe�ʾ4j��ӊ ƀj�cY��-�r.�&���>h�;d�ߗ�5.ŝJd�^
�U��E��#K, GA�*31f�-�4�j*��>
ijz���
9o�R�^zK3_�}����S��ߠ��V�z���Y:=!�� �v*��M�Mڹ�X�,TR�ж\�&��V7Ԃ��_~5��mr���̐C����������i�Ƀ?�ˡ�t�$��@ӌ^
9� �r�7��Pv��cR֒	�ᚘ��B[�8��(c��̤�o���UQ
�-�fL���C�e���F���]:с��Yd��]sb�F���lQ{�u�֮��Fύ�rKv5�&�}�p$T����Y��O�`�aX}�i���%��ERtpE! ��L�R��Ϣ$_��X$nI4�k������p�<e�``By	&KWQ �
Ϥ-�^�^4����Sy�F,��ݴw�: ���}\���_I�@W�TjC�[[��w�Д����U����A�;�ת@dL\��n�l ��{�T��AD�x�~r�g��f�]9F��	0�!��:�B�]m'�'ټ��n���G�&���q(���	1|#��ߋ����3�|�5��3�D8�$8 OO�T����Y^���t�p���ޜ*�fO��I�߯NioԾ�|o2�u����/��ޙ��r)o�>h��?ji�2~��nC9"�g7����*���$(D7�@�����7�"�Z�&�d��#Ha,Z?��x��$�>EX�U��9�ý���pb��@"c#�������s�h�'�������5w��� 2>�z{ڍ$co�Ű����`�]r��͈; ���P_8j'�e짊��q�Pl��?Y��'��*�(��1mie$�o��J��:�3���Vx��!�&Lj;O?�ȭ�`��:�ȶ'=3%W-!;�S�:�߁���ծ���&����׻�iP*w9����!��>�ҹ���Q%q�i� ߃��_ECr��KI�8���뻋��	���`�������Q����e��Yp���bX�R3���x������^ ���:�Y(@��X�_^��66�����$�vOe�HA�_���Q�{���J��߾�E<q���f��M�YŒ��,Hfd��b!�{gŔ3�2|(��������`��|��`w��Y;:y=��l��A
��T;s�a� �L���hJ�*a*���ֽ.�u��I��;D��
E=�׬/��|]_�d9��n���[��h��Х�RX�8�R�Bo�'�#g�Q�Z�V�Ij��S�����aq2��._����:��X(��$Xp��I����������{�aÿM�p
�|�x��g��^����W�L�w?P�H�Į����n�]lwl;9Y��l����滛부S5����L���F�=�w��q�5Ps�_+�101�1�L%cV���6��8ݸ��\�:���R����nަ� nݯy�I���t�?����mo����5�5�r�S�o�y���	���5�
��ǣ'K'@��6��d�r��^�3��0ټ~�܌���#�v�l$+�����Z�tQ�Ύ��W�1�*���F��@L��~)C/q[�W����T�ʐh�ϓ&R<&ԏ�!D��K��(�l��	�VH��w�����y.���Jf��V-��{�۠�
�� �ϊ;�Y��ɀ���(�(-��ば����Y=����0������a����c��h����Q�&��-�=��x�vw-[ѻ47J�]��@a� �B�:�J�^ 2�e�k�{ �>�~��L�'ʂ�Z5#�Ŝ��,��vh�;�m�qmK����y��mW;�9�+ٗ�����&`�(�5�F����"��|�}��OҪ���	k�~��o2U[S��$�V��zPl?�����ҽO�#���|�T0T��i^�w5d��k,���G�%%DG��A��G�5���e�����;W��-�%����V�P���X�?g��s2�6Ѫ����y~ll�G��_*��fp���x���6Q�"pu�W�$�[J���;��r��ċ��㲿�'W�6~9����>r���h�Wa I{�`�,�
���K��D)|���D�C�?\��I�����^V>e"X�Q���<�����',h��,!x���G�����p��8ִ^I�7�����/���%r�zKsF��/Ɋ�Q-��@��xh�u�m�|�[=J{59��o���Ⱦ h :��.���{رUr8@D[�'��E�!������D�p�����.���&�.v{�ge����l�H�M�+ :<F�k����xW���O�m�*�
[qcG8�dHr�nS鴾�C�&�� q��I9����%�j�lGw�M���x�E������Ss�;ަ�=��d@nuC�N���o�-�ˀ�Ї�:��߽f�V[.*��6�d1��JBM�e;4�b��{%�=7��C�r�	,Wf��jM?%�$����_4�[�F."%ի���@�V{.4u߲����D�K�]Oߨ�j�^��,nk�/�m.9��a���t]?����{8o��*������$J�Mɪ/�Y,�Z%���˪])qҽE��w�I�Z�ƇrU��Uy������/�X3�EV�=�����+�$�x+�.I���8�t]탟[
�c���4)/�M�L�>�c�5sH����2_v�<�#�5��G0��Q�R�����r\�<��9s���^#)Y��Wr�l�F���ה-�v����#kf0��]_��=��q����o�&l�R�6���-�p9�rf�n�*�q�]��|G�Ã�m�6`D¡� ����~#f#d��3�U�Dt@�v_1�¢�j�+y���\Inq�F5�qA����A(f�����1-�XH�i�P��^�5(�)����0��������2U�o���m��:�o��0Mm�
����<��ue?R'�����%�(E��66a�uGl
6J5{<D+?H"O{b���W͋��?�09��O�q}{�$�t�79{�΢��
�:]�W//�À�v��I�B%9��nIJ�<�;;+�ʅ[�R��_��J��776(��_'t�c�"��޳3-\}uT̟BZ\�\u�'���ܤ�-����o�4&��ge���V�y�;��Y	�x��ۦ V=#�A����B�&�X��a=��5�W��5tY\K�a6g���j�q�
g�R�~��JN�� ����£��� z�6lw?��v;�
�!���g�m$������ Ԯ�*�豆ې�Ux]=�SC�
�\�HD�M�e5A�a��d٧u�>�l��Y��e�E��#h�����������'U�n����k#fm��*l���^s�1������ o7xx�7[Vb3y+VU�4HU���\���L֍��q"��J�8D�z_�<fI�N�}�����4�U�d(��1��W�2�EM���U<#���·J����Ab�R��;����Pm;��#�el�L/1č��e����� �`ޛ�����rH2�K���3W��&E:uf�@�� X��k�|�٦Ƽ�nۨt�Ų�b3��D�3r��"w��}#�4��4+�xa������t�ޜ4!FQ�Lg�Cu���B/k˛5N�i��7��d3{��kؿ�3������C�i��\��q=��7E4��_��Xj��Ԍ1�Fj�*�Ì�rc�ۡ�b�]��]�F�g�k��z�hO:˘�`�"�Z䍓��@_W��T�k޸�f�I)����UGZJ �}�Y���ߍo�7�s��d�BZ�#>��G��1��ŋ���Kn��W����yۃeOW�b��u^�����5x�D�Q^7����C��(���V�,��adK��ic�k��#8��
���x."�[bcf��e�e����u7
WYJ��;��×b�l~|��Jl�ؼ��wu���/st��!y�Z���oN�~�"�ZJ�S�Us��᫪�C�VB}|��<t}�.�'��!F�ɘ�V(�fi����)R�mr�">?M��4k�I ��!^������W�}�7����O^\[֞�_�7�O@e���DI	����ǘ�H��~����%��r��r�Z��?�o��9i�����׳�l��;���v�2(����x7ָ;$4��'�����M�<��qwMpk�=xp��;�Ss?�יzO�/�j��o�:g��9���%>7{��Y[���W��6��M���[��>"'��A:èC�X?�H���	�a��u-~��B(uh�%�8��Rܰ<�Z�X�����~%FV�t�M�*�щ0�z��:��횼D�d����M���Vy	7rd��j���kÅ&�SKj�P�����7�5Ȟl��vK�X��/�+?i����O0UE�c����kV�̬V� !�XG���@gX@ۑ�PV3�A�ք��nƂ�X�qM�F��Qv4�)|x�z�bw~P���]�֓�o�u�+5�0Q�v� ڦ˪��/B5"�Q����ڦ�r�6�+Ѕ��1��g��L�6�T�"��1*H����aTWU:`��%�Շ����3�����&[>�f<++pFb���DT�ȥ�hp�3SR �7Q�Gv`�����qg���A��)���F��ԯ�ۀǎ�V�p����f�L�4���ދ2��yZ��LXh���o�S��] �ߕC�dy�Œ�dVJV�Z�bү�\�v�0cM.�&^�\W����s>��칈]���He���:p"fh���+���x��c�J�	�O����ы�T��[�I`����u!Yu���}��M�d2%L	�Z2~�A�֘�)	Bp�x�r�� c՜pZ������|I<,��8�C���0%Z[̈��Cر�T���C�����Tҳ%��	����`;�V�խ萳X��-�5{�*P"Cx�r�_y�%j��3�B�e�.]�`�?�M��9\L']�Z��G@O/;�[3㴙�E��^�g�K\�W�>���MEk�2e����2u�t��p��D^Y�?-%A<iй/���8V)_�l���/���`�-]�����MG����k�L�xDŶ�Rh�۫E����I�e6R?gb�*P�I_�
��F�*��烻g�(���>�½DBy�C�gZ�~�����ef�y��br����d����zҩ|Q���ׂ7}F�B�������Q֌;0b��w�Ws&�t@���11�B�󋝣�Ж97.�����aæJ ~�&��7������>˳��\(�a��T� ��������@{��ϡe�E�Í��M>y!vhcٗN��dN$$�D�lr�. ����Y=5H�Z��[b��]۾3O���7�������4��DЍ�E.�'�V�du!�]�����z�M["ߞ�HfD�cD�pH�(ayP�̔p�����"��%��>)�sbZSHB�m�6��T�qB�o�D��ǲwD-�F(^��F�v�<f&�#��ם�����.2I�bST�؇ә��"M��>:�1�������O�pe`�	�~F�]�W���[ �����Wq	Z�4v'�BuFV�"a�!qz��QN(�iEx-�Kc?�7�X�ׅ�e��m#�4��tĚ�X0wȌ��^ �:Hj�VH�"�(eF��ڐye&�{cX
:�\���<�*�c(�"�U��ւ����˪�+_�G!��  q��rgH�e�PsX�9���kՒ����FzQ~�{8ޔ�^Y.��>��gO�˼�m��� )<�M9Lv��{Eѫ����r0��kNܘ��Q���]hﴣ�U�:G��>��U�&a�gXH�S���;�}X��F���g��9��ఴ���un��"'�i��h��<_Z������{�@�r��a����7��ryq��κN�z��������e���Գ��!M��w�m�S�e�����r�z(�Z�ギ�b�8'/DM{�"o�[*[v��1�J�Z}����
�)�MMt�*�WvV{�q���:tMn��C>i%�xt��;:�`�vN0h��ަ8LZ��<�zƻ�ps���Z����������g�FfN�P�mz�����޷a�g-N:��EqP3���vvPH�]�F�5aN;]��Nyf��rh=�"w{��>�秅���a�Rb����-I3�Ro/� ��\��\���Tl�%/���̻�C��Ab��lB��Bw߰9�����}6.Y�� u�>q�;Yr�h`x�G�|�t�iO���wx4o9̴�b�I #�Z�@�*B]w����}XUd�yӪ	�G ��a�+�we�R��k�$�\�g��'"�t��׍Ҍ�Ƽ��!ԁGx�A"��	�Lw>"W#��7�b[��G��>S��)�(3����)az/4%�Q�T����(��/㔲ښ�!{��6X3�x���v[�]���/|�F�❕\ԃ��<���=�K��s�����
���V�t�.�u"�S:���xw\��"DYrB�>psi1��4�W�{�*����X�3���`��p�������c~�so��N{��cծ�aL������R��{A0]��������kk�~�����n���C��߭4���ь��d�>o:}���`�]b}5�^�:Q3ăM��e�0�@�ϸ�P�C/赋�:!�_�t4���(=H��,�a8̰(�=����s�3��Y�^^�G\�Q+f�n��;Ӡ^�K^��i�6��L�����運�?O��ۊ��u�h�	S�E�w%� ٙyD{՘���X���_���)�"	�d�5&2߉�����0;Յ��O�� �>Ғ���x�#!ֹ��`�އ+��)X�t�ﱼ��.�p8���L������1Fn��җ:>p
8��RW :���wC<��i��(4-n0��~\�a*�u�����a5�Pb��ڮf*BY��5ig\fhC+��c��0�4��C�$����q!cvp״K�`NxW��5Z��+,��2�/.Ī���=I���.�A����>��T�;#�s���~�����Eu��5^�L�Q��Z�0�c �?]�#��GE��$Ċ�$�r�ِ^j�Oz���j:�v�Za����cLV} 4�k=�|�I�����w3Iɉ��[����=�:JMxZmM�M�@�'�N���_�|O(����*|) Q�?�9?mr���5("o~�W��b8���ϩ��Ͼ�8�Iii���-r;QV2�:����L�,��O�Gs�h�zas��M�)S!��MZ�=��'9��b�}!L�s��P߾r���Rǳ��N���0z85,f~�"0z���ݲ�ֱ�o�2^{�qk,8ɍk�}�Ra��y���Ћh� �\C��@�~�KK�[��Qx����/.X�}��X Մ��aF�����R�sqh*ǡ�PB��R�C~�-�$�e7=;a�Y�w��H7	�o�/��DhE�l��J�|ђ?�NM�/qr��5�1����]f�����!#A[�wl��╟�����F7-�W�u�0 _r���y}7 M�o��z!F���ܰ�Ym��1�8�ڤ��Q=�	/�t�E�v�����W���p/�&5X�G�[tI�NΖ��i�y\r���_����W/�!��L{/?\�ȩ�e0�,-�ۭ5�*GL�����=v�=V��j~p6��i�V��µ#sߜ��3��3�
$^�|9�n`�f�X�NY�������GW��|�z��Vd�-Ig��gvݢt�O��ѣN�Q�iHC��q����,��q�z��9��d5-�����ϻ*���M��p��a����<]���#��4.��!;���%�%H���0+���7��k�d�Z\S.�UP���|/xl�`�����ߣw�HL���Xf�+V"��Q��cm�4���V��na��#tj�5 g{��t�C�ߥ������#Ǧ���#��U���4ak!�Z�Dr�O��\�q��x�AT1�}��geL�����g�?#�q/0�20���"�w�49>�/�g�T��:M��p�e������WG��(N�S<�h����iϿw����eyC(���-T�{��\�����r�F`���}�?��6=J�?+�ԲagX�qq*s�z��IM��Ԭx[Nh<@����� ��5��}N-���Ŀ@<�$;"�����Y>���ꮗ|/�̿��p]Uա�g�ȣ��H����Z ��9#�k[�,~	߲^� t�����T�-����M�׍�����v����N�Q �� �q�[�	ge7*Z$L���\��w���:�촦8`tL/��B�}k�[>���YR��T�FŹ�G�#����v�N�!�A�Z����6s1sLS��7���������n����_�ⶉ�wԪ�|�z#�u��=T%�У_1��+u��ŧ+�*�	��3��2?%".(!kk���M�k|g3i�9�4��8�~��?����y9O�m v��`��ֺ��(�2#p=����|�)��)��+�B�j���e�[Xd��vǮ�oZ� L��$�R�x�{���K��t-'�A[/7�!~t�īZM���iD��Uu�$#��ӆ��,�يi�Z�ĪP�v�zW_N/o t'e�a�=�q��d�s����4/�&T�!�ڏY����N+����'��>��|��bqEg'&"�1�J��?�os'��<������=���l�	e[.>��;�NI|'*C��tF��8��(:k�A�kx�<����箷� �#��lJ�K��b�
��Y�[�xY�á����5޾�#�a<�*@{��f�~�@)�����v�攱���=ܯ���&Tʍ�2 �����v�Y�v��֋�Ƀ�#�
�qկ���oa�+O�F��f���T�4"����Ue?�9� 0�U�5��4�EW�'
J���j���{�����?GR�������~��i�Pd����9�FN�C0�֝j
�Z�5z�-�d˄���[�n8j����6��+�.?!��F�1ө��s��*�ӑ:����6
TP���#�pt=�l��v$�S^&�����|�J%э��R.�-`wT#�ha�#`���ݬ���#9��\Q�1��u�x_�m`#�;�*2F��@77d���XZ��p#v'��4o�Qâx*�z]��H����iR�����	�Z�ѿ?
��{`cMؼ8o\�a[o���:�¸>��K�Z	���zqN1u��;%��
=����/����H���bY Ģ2�}��j���y�a��X�#��n��i��ËF��]@O4�)�r���C���D@�c{m�A�r�>n�z �9�h���ƭӑ�UH.%�k�)J��j��U������Io�i�6���#cC�/ٜ(�;j�+]��r=*ݴR��!�;�gc�lQG�`
��o��jKs� ���$��ꋭ��}|��rLk�;.������M��
h��Xq8e$�z�A�rs��.���T��X�1w�9�HXo�D�J�s�0JM��whK��t^��Ș��Ѷ�t��W���R���W��d���-y�%o��?;�䍾Qζ�V�R[��d��`)X�rE<�����rt� �Wl���$��!S2o��7����<�;�v��̓�h��¹���ϐ/��<?%k�}{[��沓���PƮ��?���~�ٳ��m+�$�a�hXڬ%��n����<]-~��D���I4��bD���.��
MdH�6�%)���	�k�Vh��Q��M�bU�y֗�}���3�(�mo4��i���D��~kVU�e�����غ]�`�~��6���qn��?݂l��b
p��ܯ�i
�>��\��:����y�Z�Rz�J%��Q"Uz��XP��k��{��Id����Rf�ઢH��^Q�j.��<C3#������R���֩81������=O��5ҍ�m����u��}/O:I6R +�H�aۙ��*�@�H�h�����M5U�L�Cr�M��T�V�Z�ٯ��\���s�gAx��, �[|�Ҕ�֊@8�a�����t$�kیֲ��Fa�h{> ���֍�4�IͲ�m�]�7[nI��)��8�Ľ��093��U<�����_3/ ��J�i�A5\;���ͽ�\.�w��c�h�¼?�=��-{��iO)�\ս��|q�"L��-c�8�Y������ݛ�J*����hG6��F��z8ҩ6��~CP��k
���k�\忡S
�{������R3�9����#�/Ҽą�+}x)J%�č8kwt���M�7>����P�������ꋟ�WOb�ǙQ��"r�)lB�c��t��ǖ�S��m硙��m��f�	��C�Vl��GC�K���h���pQ�`���6uT��;?��n4�������W��O�fZ�����m�O���
k��/�a���\���.���!��1q�J��%C�����S�O�&������C�Yщ��7p��+E��z��A��E���i�l����)/g\�38�����r�I�,ĝ��:n>fbb��cE��#�=����_��t�n\�Uh�R۔��pt��^)���&9�=�k������D~��ش�xUH�ݣ�F�Z��,I�Cڶ[�Y�Go�4���R��� ���+Lu;}�I
-s�� ��B3�3tg�=m��x�\�p�����,�͎oh�cV}H�lƥ��r�eI�%�J0�r�JjI��A���;箑����|�Zݜ�g[H*V���إ_5`3<�^��MuG��
Eq}�����6([�P�#�Θ��I�5#�ɚyP7P�3 ��@��\
�vci�t�F���C(ï�ކ�G�~��D`�t���� o6{��_�����\l�60�W�t�?�I�K�A�1��s�x���O;"6̽��%���ˤ�dy���QQM�:��n�]Rs�A��R�n!�98[�y�~S&eUv�Lr��~C�n«F�)'��8�o̻�����Z���Y��}��գ���Lc��S���qhv��Dcn~�������D�\��}�X�@c�r��^�m�{��?�V��噅���!���\�O���|��N����j�=���9d���<���+�̴T]���|�8�;fh�j1�]��DOa�J�|��I�>�1lb�O,H�:$\�D������m b�iy�GK~h�ظ)���rbE)j^���Aw� o�E-\�ۙ׃���2)Y軸��1}&��eʥ��５�*dq�>r��+�ly-�'�%t����Wny޻G#��qF�/�
�3ͱP�M�F��w�9U��'J^��}��r����v;Qi'�Q�����z���L׊����9b7t�*1z'8d����D)�i�Aq�|#[��Q�x���P�v�ݸ5Τ���_�\�'�ʱ��u/��o�%5���� �����;`�u�m���m^�Z�)t���H0�S�Y:�`�yWrg~-��+�J���+�|����y}����яb�:9j_��hn�d��+"Ci$�PkqC��agv�Z�@��0����̛��#���'�:y	39���$�U'���ɍB
3j��+�q�I˪*䌏@6f�a?溦�O��{w�z_)��1=u4�O�\����ǵ�N��u�ϻJ�&2(�Y��Se0O�+ʋ�V��,��
������ݡ4������c>��M�Ad�����*rヱ���c1æ<$,�Τ��z2�1�DUz��7��N��,�-��I��!ZBμ�i�����&�S�/]1$��s�ا�l����Ы��3�>�M5�J&-�%�����2?��t�ǘBjQ妟gf�;W��Át����V� ��௼nV�qi^p��^�P���<E�vW:��L]�}G8���W�*�����J!�y�����%u=;���ϑ����7,��VG�B���R/�ד�Q��RUR���[��#���	���8O��!��1C�<vwt��v�����1U�m�$l�jX��-�%Q6=<VP(�<��7�*o�̪���On˅s��7˟T�0��2���p�x�ߐZ�d%~��"liiY�9Z���P�C�@NvmN\�Ir	�n�� ��͍��fӫ�R�j�V�%R+=(��N�i��Q].q�Щ�K5�	�����Z��tG�����)��˶t�4�\O6�	l7Bk�h)���*���.*�I
N2�k7!��Ge�Z��ԡ=܃r*���-[�5��b]~,�E�s&D�}e�a���N�[6��;�4	>\����k���=6�2/b�n�Z�r��f���ITP�u�d8�6oXD�,i�j?2����0�l�SM�D��$~�=b7l�A�������*�Q��J}86����8XD���/�~;��e=x�^�Uwp�fք�!{Ϛ��x�Yl��b����X��	K"�j�E=��~��	ω�3y��_?]쭟^h�G��QC��IC�aFu�u��Id���׷އ�����ab���p��moM���Qw7=�"�^�D�3��`r����g3�-c����Ȟ��\i+�7Cp�D)ݘR:�~��b��N�1�����'�H�2~������,1p���w#��!>M�Ʌ@�o7L'C�$P>4П��>z78���F��>�5�0�	*�퐷�p�&g>#q��F>�SQí�^���\��|��|����lsT��]'�����v��W?m�����E��v܍:�������}}
��݇��Xg?�Z��?�<��UP=�#�x1j�JE�W����!�(�Z��ax$I1\����dU�q)�麕��0�2�=^��aB$}������<d�Y�������o
v�t0�l����E��c�U�.0�M��~^�^	�W�5V�{vc���_���0a�M��xq:�F�)�_"3J.�/|i�y�y����~E�;X��K�$�
��daL�cƫ&�ʷ|O(����Ʉ�P&���l����l���w	�
Q�5h7y���S6�'�%�Y]�O[/����Om:?W\�5AV�{�i����"�~C��Eq,�<3^iJ�v�M�����\%���L�"�n�5�{jnaf'���L�=u$N+K0t ��*|h�2f�G?�9�$�ӅWS c�����R�&| 6�]���c&��	�U��G��p5i��.	5e�9*���PVkf��p3۾2:�	3��,J���c��Ț��n*���嘒��͐�1��aކz�]%H��q�37�:@�v�<�m�9������*W�'�=�{�gs�IZ,���>9�^@�߯��^�+�Γp�0CXn�I������B�[�#�q���O�����ץ0��ٮ=�y��<_d��uݯ���t����>�^_<P�e?^����#�P��K3Q��2`z�A��7�8an��`-o�j�a�N���~wB|�7�P��Z	8�!���/���{�;��շ�B-�V�׻y��x�<5��������*D���C����Wt��P�`񻴡07=�pn���H��ܝ���ÔC�w�1:����Aڼ��-F���o�7u`��I�^�_�j����ݪ�&��B~T�=���C���*P`��av ��J��a[���VJ�e��V���a1�{  �B��w�U���Lo�����Y,��f�X��NJ�#猞&��}Ч�&#�k�C�Ͼ��g6�G��ބ�S;R΀=����e���[D�ǹ{*��"rؐ~�n�8B�T_�-b����:��3[��Q*�|�E��li�(��}.���U��o�@/�m��*&����&&�-N�.;�Y�w;>��
��vL��@K=9���	1�סchV���-�6������we�,&��~���K��<:F"3���Q��]u��	<��C>��h�����f ����x(��[4[�5�$���՟&6�G�&����;���ª�/�TQ;9�X>R�B����!)r��^��ђ�����7C���]z��R��i���i�\�
�{�B.�N�_:r�ˣGӄ��
���xR���cF�'T�CQm-ck��GyY�xN��+�.)S�oCƦ��u��Β�hEgmǫP��L�s�����]�,3�d�`=x�����5,d� ��7�i߄�f��νϵ��An4�2_��s�T�R+x|_Bp�D�g�B���!6�G΢ou�'�R���w�B����ԙ��z���:7�Q�5�]�K�Y�w����'�l_��bj�O��"�t�vj�_�L��ڟz���+�M��cK��.z��A}.��ߔ�� o�6����J�娽�&Ȝ����D8]�+◤����O�KS챔�^%|�U
ִ�PDs�vw�)�����ל˿��
��ZM��E��:�2�`/g|�#�WRS3"盚5�%�<n'T���欑:�y˩F%�\�%w��M�wԃ:�j��Tmt��������67Y�&��G8��X�!OW�1�E�W�r,�Ge�C}8�l�Xb)����z�D)�$ lqښ��a�M�%�#}��h6c�,̀yD� �⋫f�W:�*��ڂ�}���ŀ���K��C?���GT,*2f��!���7f�o��B_���FWҥ��?G&����}O�G�����zqL���&��P�O�����7��C%Yr캒o�o�����:ϔn��64q�K:]�E }���9_]�Q0{D��@�w��NCq.\��TGNŬ	��Җ-�~]�5H3mq�O�@��t:Kl�f7����A�A����~�g|X�oxk+]!�����I�Ir%D� 8�8�V)i�ri΍������<H-ĸw�h(���U�$��?B��ÏY4/��������]��d�ϑj��94�n����i�*Y�~*�����«S�ė�&ASx�e�Ã�'XY��.-��n��+&�+�ى6����}Q���|>=�I�W����7���w'��IR�JsΘ�T!�2z�(��"���7zDXT{U�Či^!jyy����`_�_�L�ib#M��2Ԇ��&sYE'���9��d���c�Kk��Q�*8���{���,M�u��W�)U��i6U�S�����_��5�:��삄7�f� _�[\
}㞟�On�O�O
^+���tl�����!��n�]����!�uP�ܶ��?�<��{o@I�ò����^��d�q��dŬm��=n^P���d���;��G��8�p���h���-K��� ��Թ����L��T(��G��F��b�!�22>1,�wCƉ�����v�N��ܝ-#�"�߶�c��/��h�en�8�J+=���D=�?]�H�n8oԥp�	�����y��CN�_���8zZ�9��p��"����L�j_��uĿA 	%t��B1��7aZZ�S|����c����oj���&��Wſ�gAA(+!fp�łT���F��5Ǘ#��O����������?p���	��
2��������_�=�E���M�C�{}�Q���4��/PK   lV9ZD�h  �     jsons/user_defined.json�]k�0����-I�iӻ1o����2b�j�&]�ND��;��`�����ғ�>ys8���F�u^��*m�DzS�kk� '8!P��,�zT>o?�|�N�|=XZ��j൙�G,�1��୚[�!z�[�[���<+��TH9�1�B�E�	�`8���e�:u�4V^8ݴ{ß^�8�4f�F���,*7�t˱�<����h�fI�sʠ���ޮ��b?����,��|h%�24X���]C%��唐��KH:�4ie��:��Z�

��~��>8�^�ڟBO���\z��N(>��L���lF�x|���n}��\i������r��E/dFX����/��D������PK
   lV9Z���  z                  cirkitFile.jsonPK
   ��8Z�=�:��  � /               images/a3896090-6cd9-4aa0-adce-88a16a68907f.pngPK
   lV9ZD�h  �               � jsons/user_defined.jsonPK      �   �   