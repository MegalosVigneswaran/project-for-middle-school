PK   o�5Z��N�  �<    cirkitFile.json�]�r�6�~��rk��3�Mv��Tm6S;e/f�\<fT�H^Y�$��w_��e�$ȏjHr&3�m4��C�4���_��m�\�������r1�a�j�>]����W����v���i�޿���^���/�|��~�(�[��T([E��U$��QZ$,b"W���,��m<�y�����V�ӪZu��Uֱ�b"��<�d�()�2b1���,,��[&g�=c�	uy]k��e�Ge\&��3%q����$�F�J3�/a�m�5i�a�bB]���َ)�mh�mi��Z���^aD���Ib}�Zc�X��>F�K<�"5��&͢D�2��(�,�d,sE�HlI�r<�u-�Ҙ�W�u��"J�P�b��DQf�,g��m�K�<Ҏ.��*"[%��یgU�Ǚ�(]s_׈��uM\kܷ�'��V9�d�u��4�"��8g�-Ka�N�S��K��4�{�RD27q�hn"S�Yi���)�]��SA��P�V��-�Aڐ�O'a}��-|J	뛴>�O+a}��-߰���9��q�����:�dbt�1�Ee!bQTJTI�=������X��Y)+y$�̣��eT	��X+�r�i��~������Ĭ��s���$Q���u������M6((׾�&�`pȄ��g�@A���i��LX����k�|a�M:����N|��Kٴp��4w���*S؂�L��{'��<�Yn#�3W����%��<�bEjc�l���l�k�d����z$>�i׾�'�d%����6�g/�(v%�Ҙ)�&p�/p�I ߡ /]/n�Е�d�4��e	�2�j�;٠ۮ����������\��s�6��I<��|
"W6�k�u A�� p�2�g��mЎ#x�Nq愸&�}��ٻ�)Hp��{�L�+\�$���W��I�����6��g����x-�g������YPz���y�O/h�Cu��������T������Ũg�2�I�����3O�[��.�3O雤�i���#-q�\>�._�˻�x�j�u�����AZ�AZAZ�u+UElE�Ei�i�i%	��@��^�,~��L�0fa0��mQ̔�\уo��fTU�f�4�T��i��F�eM��A1ߢ����%|If��N-פ�iP̍���L�⪴	mn�FR��5Ӡ85�HҮ۠X�L�6�ŉ�iiI�����(�Q��i��c0�z_`�4~?�(�X�/`l|�4T=�:V�hx�4,;�%��x�h�rd^�h�0/hpolMc��a~o�h kxDh`ixDh�gxDh�exDhdxDhLc�l��'Fd�Fd��G��ӇG��ƇG����"Ǝ���9����s&��˨冺��2�}����o��;|��ݸ��o�#;|����Ӂ������N�%��(׫������"��"��������b��b����A] ��A/_�,�Y�0fa0���A1�bH�A1�b�<�y�0(�aP�àX�A�E1����2�����2�����2�����2�����2�����2�����2>/�ӓ�
��A�'��0��nذӓ���`��`+�ӓ���`���NOz+�2B�����NOz+�#����VFϽ�ӓ���vz�[=��NOz+�'^����0��>�N� ̈́����ӕ��������uv�����|U>��ߥyY����UQ�f7o��E���O'��&~5HysH2�=]S�)�OK��5�_�/�(��G#y�(]S�v�?��5~��y<��"x��a~�2pΉ�~��5����I��璂�O� '����<m��(x�-8�%ɣN7�kC�b�I�l.�`�	vJ�H�K���J�S�(���b-�RK�Y��&Pmʑ�y��ZЂ��Y3�{ΊL%�b���צ6JR)�J�"��Ƽy�����)�b��&e��o�O�~�QS.���!ERI}�f�B]b�0�Ag�)�M��K�S��\��;�g�.ճ׏p����\'��]�o�����O
��s�-�O)!ϋ�<����m��qr���"gd�ܨ�=^V��/eq�.�� ����"1���I2t�q�A����Q:�`�b�f���9 Fp�9��#�3��9�:��#�3���<��#�3��>�3<g��З!1 D_��8��p�Ĩ� g	ї5FDׅT���P#F'ے������#:�0����a��d����P9�$���!�_*tK�s��!�+qpU@�ߗq�%�_�T#!8���CO��]C��+�r�U�����w>�bY��b�7���\<�A�8�^C��6B Nj2��n��:ԛ
�����⽅�20�K?�-�ǔ.��'��j����x���n��c�Y�=\؍$�C�A5�h��G�g�»�Y�*�]J���˪�4_�|��l����sb}A�_?k��Qd����.;�ϢPر��	]dxR�ɨ eT�6/�IPA���#5@�!�����ZW�����\��H�%�G:"SQ�{�'҂' l����� [� I���I���	��Aslu�K�]>��?���S0��1��Ԃwp�A�;8�`�5J�uwh�A�;8!����՚GK��	1���wp�B�;8ia�5�'[��C�b���1��Ć��(x��	��,��,��,�,�,��՜/r�&H%�fJ%��L��N�'Q�gS؜���p~ŀs׵.|�w8��z�s-R���p~EJ}�c��v=ց�z�s-����h<�b�=�ba��O��Y.��f��̋ڻ�:x��ˈ�V��^s5c�����\/�zi������76��fJ�yn�� �Yf�&`5=�+��F���M�u��`sO��5x]������j�P����;�M�̾���Y��`�T@샃
ȑ��r�>�8ض�u�px#W	9du*!��nO��ߩ��L�:y�z��q}J[F���fyQS��(U.b��	ˤ}�F�Mc��L�&+��bK)RÄW$
�aRE��?b�%y�$SzC)m�uR�(�n�2u�HTf#	���U%نQ���;�J7dQ�kr�a��sn���=å�⥜q(&�N��P�N�Ų��{(�ſI�>R��U�<����HG,�mD�6P�Y��Oqu��=R�\ �dT�3�tmx�H�(i��<]"a�=����D{FB��Cy��g��F�GB�_Fy拧��Ɣ�GB��Gy/��5����#9S^®��9Ua׳Ba�����8��CNh���!�8��P	�P<[}���wiV���_Ko�����jQ�Jض�u����w�ԶHu��Hv���Hw�̶�t���v�؎�.��{�e�q6e�[��?��=�u�͞�~pRI��n�U��2]��������a]�E�[��D	�N�fZF���l�I�2�n�����z,����]Y��T�����M׵���O�V��r����S�����_�6���z5_��F�H?ԿץW�_һ�������W�0������u3s?=�_~�a�kyvS�w�+|(W?���]��۪���|U��������J���Nj�ga�왗oV˴p�	�J�����|=_��x	_�M��d��*�B_��<�I����ε1��0�,���+*�p?�z��s�eE�y��拇u��7u g��l��;���f���O�|�ߕ[��ܚ�[n����I�+G(�#Tr��]�������c1_�X�6}�k~]{��`��dg��G0$YC�"�@�Oy&��V�g�"�A����L)X)�\�4ʄ���&�S&J���YeL<P��4��`K��G4�Q_ s���*{
� Q3hﲇz�
��e����y�Cʨ��QԽ

�"�Q�_7DոP��T��"�@�g]��L9*��8λ_u}h]6�M���!�������u�1�t%��f�#������dx�C7\ ���/�*���M�X������t���=.�˟�#�U,�����ܪ����2�<���DV�(���iYF\���8�U�X�e��� �:{	u��O����m&m���̪p�n�!�����YŽ�m�y	���T(���/��t�Bt�@��ۮ��O���}�i �`��)�`7J�. /��ztX���Khb�І�Ŝ8>������Y��ʢ����WN~�,��A���.]�׿�u��Ӯ���l{�Cq��9��jV���}�ݽ�����߿���Tr�di��O����vy�܇�33m��]5���\���4?y_'OT�n����������=�7�Z.֯��-{[����L��-����ѭ��W�,?�w��ױV�ibi�rJ@�ɵMO��%.RY�eƣԝ�#g��H�V8öJSY;��c=!W�ǵ���俜i�e5�iW���j����٬F	øJ��ף�v�SņI�$�P�#� 奭ǻ����|����F�ٵ[#��*�n't'dc�cf�:5n���9Bo�^�b�;���o��$��KR_pI:[�Z+�p���'͚t�U�$�ml\�O��s�-�)~��4֪~^��l��wR8�(���b-ǐ��2�Ȕ�Ed��##�<J��fQ&�_�2���*^�-;t����^�MH�����K�WR_5y��엨��_�;ފm	O��p�W���U���O&ZdfW�k�J��u�ʭ��7��Se����2�엹�v�7}P�ʺS�+b�nj�+�����E��ߺ�+R�ݙ�u��):�"p'�����Z=��_}�(�:n ������1�y�Na�j\)c��ˁ�2�Թ��L�62�Qeben�kec�Y�}	���TC���C�*5�L����C��r�L?a�q�i�VO1���;����z��$�Z�W���t`Y�j�7��`t�o�1�е���=�Z����O���]eҥS-�����٨��ҭ�Y��=|Mf������['���|�~_7�j�����r����԰�ڿ���vؾ[�y��/�ovoD^�����������ߞ��֩?wp};�y�td};�z��N�r��wESttփ��rQ6�=to�Z�_�d͵��p��/��J�~���~��C��.x�����7o���Dn[�����`cd�>��}r��JD�˵0A�8k�8'p7Q��#�l��_�8��Π�<����y�ŉ�ԁ�	f���9�7@�S؛(ύ��,*�Y�m2-c��6J���#�d�M���q��:^�L/�"y�� 4���&?7��^��p�M3,��	�]f-��:��
�sa�N�cck 6&p7�avO����7t�Iw
�`�
/�	�] ��  �?@�d�@�	 � �	�MҦ�	�(0 ˴�d�@�2�5 8wSr�g���O�(�F��� �e��@&pwi�ȶW�;	@�<ϗ��e�� ҡ���u})�L��� i�Cw
�L�y� ӂ��x���;�}@�(��� ,Qz�p!�g�sG��;<;��YqB����g-T0�(q����0Ig��pq_�A�y�Չ��,��
G�`~踗D�9����5�E$Zd��n���Q����^�.N!�_/l/k\�y�.3�T�������
�aT/h�L�smw�����|'�q+��,k��p��	�jk���G骎��/qt�� �?4N%��{8,�	�M�	Z#7P;t�����V �yp47����d���`�}m.���hwD3�@xq�_���¤��`�����E�Zt\����|G�y�4
7������F����FEXu����S�흠||�t���S���tppm@�oj^!Sx�,D����i�yHG�(UU:!�}$B��T!Xu��H�:�M�=t�H�S ��-�C&I4�Y%�5�#�	h´��\�kA	�÷Sd
��yb!�׊q�L` ���{!:�C�9_<}�l2�) ~GC�$���!�kt{�!��CZt���(�t Dtj�FMb�����N8��	���Iz$@$�C�t��������N��B�I4�Q(D&�7"-��W����ѣP�f?Dm�D�������1"`52��� �I�N�?�VG��Zi26#0c�@hϫ���)�MF���":�{�h�TA2!i��3l�s�a���>�)�MFH{��Ҧ3����d�-�D��ڀ	��a�\0��j�kP���l\&>�EHi��1�:'֖�P 9.'��Nu����P������a��ɅBRy��BG�QP{��ޣE �un�������\�ӻ��M�������t��}���ݺ��P��ݧ٧�PK
   o�5Z��N�  �<                  cirkitFile.jsonPK      =       