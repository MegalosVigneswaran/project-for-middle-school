PK   ;7>Z[��=  4�     cirkitFile.json�]Ks�8�+S�UT�E �mgU9�&�ٚ=�.H�c�(�����M��/@)����rCv��L,4�~��&��l׋r���g�l��urE�Yrk��y�-�%w����,~k��mr������ٴ�|�۬�]��*-��RA�HM.�TZU��WeY�I�>Nuf5g\�"���HE�L��MmVJuM,#Ɠ�ٳ��nhDw��*�L����p�
[���%O����T��Vn�Ɂˬ�eA�(�u�.�4g����*R�i#���}a+�cV�c�LS�)����ROO�^�Uj��w˝�y]���X������r���#u _ �	F�Ў�Y`F�AS �.B�]RmS����dE��L��H�e�I�	nɲ��u)rF4I���W4wl2����_FQɂmI\2P�Ba[#xe���9d>��dzd�D�*��!=�/bd�5	���sȎ�F�6��V�aCZ1�jg��A 	�@P�p�	4����_��!;ܖ��C�^ F�pʒ��
�]��H�c�	r�P���a��?{	>�DE"�ǐ�cXC��Cō!�	]��.CB�!���%Bvh��y
̿#7Gn��0i�9��z�D=�P�P�-7�M�,�&ojɴ
�����>.,
�ͨs�#p9�.��Y�&�M%,��"��\rZ��@p����3�֩��Z�J�PKH]�*�1d9�]hI�,��NY���i`��8�%��4�ɀ,�rH.����)�kZ������G��q�@�	�-&�0a]d.*
�Ku�����b�q��A0�a�4�i�8(f�lp3~*+ �bH�,�Y3}*��"H�㠘�A1��b��8(�qP�㠘?E�c9aۚ�b�	k�k�B��\X.�p9��亀�	x.q�EDᒝ�.'๜�����rRG�r���u���ih9�����<�����	x.qd9�ip9�夕��\d.*
�Ku���4|i��8 �qL�@���0�b�,�Y$�,�Y�8(fqP�⠘�A1��b�<�y�P"�y�8(�qP̟��~���G�?��XV$WTΒ/��nw+�R��r��4�m������:'�ra2ᮇ�"O5/�TS�3Z��ʫ�m��i`C��Р�Ι?��ApCKT����e�[��~Э��j��4��t�I�KP4�>sE|2�MY�Q����h�ja&rX�+���G��r`d`YSXČ|�9C�D&t�/b�aꊁ��vS]��π�ُ�4�oH����4����D̺�JJ>:!_/|��$�ƎG%x�<%��t�bZ�Ʋx�!m'��M�) v���nf�уR�]�o|���Ƕ�?�-��cd�{�%�&�4�=*�K��x��Q^$�/2>��H��8���Cz��/��T�2�9:,A��x	�Z	���	_?@m�)\]�)A�Wx��,c�%�Y��E����ږ�n���-�G���|��������?�����/���`_ 0������aG��_p��[U����
٘�����w�d�K0(�o��
�6 �| �tk
�7
`�_-�D��;�MH�U�[�]�o��?���_9�!|�`�.`���0�%����F�ϱ`C���j��'�N�b�E!�bqH�@�X$2,�pb��&l%*	��a�ɰ�dX`v7k�ʭsp��� �ca˱�cqʱ8�X��=N�g�c�e�k��� ��������k5!�ݸ�,�aQ��oH�392$s�wt� �c'�c�:@^�Y�3�� ݗ[iG�)�'���{"@=uW���]}����`oߣ��2߃���`�GWO�J�������=���}�{8�7Y���Y�֣f�?��� ^K�{%%&=�Typ���
�^�̽1�4LESvC�Q��~����_���M'��_��WǏ�_Ý`g���S�j�P?��;�<.��~����������v����$���O~���i�D�M��$�M�Ф�M�Ф�M����M����M��$�M١)��Y�EcMUlL��@כ�j�m�zx�N��<w�)�j]�啹�+��ڰ�t^r��fg���be붋��Y�<��3�q�}�z�l�l�.���6�e��$�ǔq>�Z�f�a���9�����8x[�i�RS-k�*Kz��S�k�ڢ�ҙ6�G'.Dmͺ����d�,��f/S��s_�˦\��4>���yփ��Y�y873GH���@�LC8�t"��l?��j���ۏ>&t���=`�U�,�\j�˻O�4�es%)˴�'�j�p�K��T�U�
cHj��: *��9Q�P#�`��y#�dD�b���T��_��/��Y�2H��,3*z��S����p�i��{h��B%�nʙ�J|��S�\I�A�Z=U���.P*�K��t�(���ye�,s�Umz*�`�M�Ĝ{�1X�N:cG���l��	��v��n����Qn�f����km>��}�,�lV;�׿���R�K���Kg"�����˻�_��6��u�[����.��}�����-떻u��i��Y�jS���6�DxJ�(ˇ;�����:�(C�9{G�&��J΢=Z�y
4�Kf�t�����X�rcmʤ$JgɻM=��rv�$��§6�-��U1�*Uz.XN����r����u��!E��Y�l�Ҫd΍��8�oBkU�2����A
`��$�;�%�l�>N����V���/���ݲ�����>n&��e|�S�s���t>�y�OyF�>$�=k������ٻ�%d�1�R<�撪�X%T9��drȃ0�zǦ;�Po��sL�o���2J�D�L���gn�s�	��a�ʧ+�kJ�*���q�
�,��n�5-$�/�(�+���B�y<��7��ͨ��݆#��A`�Bt���2 ?Mzs�:A���8�n�m�N���!:l�t�1��f"�A�P��3Ay?r��=��z����������F؛&�}U8�A�ݑe<8�NIO����|�>��ʧ :	�'���2�ps蘃g��Y��9��{dS]X>������NY_i���U"��H��s��v�:���� ��P�˲jo=�S9�~�v��m����5���?�}������V??�;�7�m��ui����3�e���I�.������K���ٵ�#LӾ_��V]ӳRt��:�
�ܡc՘/b����=�tw��}o�ێ������W����}Ç.6��o�>���(�~]�S�&�z��o�d4'�Qo{���'Z���3�{t�i�w%�s�| �G��b9��u-�d�0�óI26��I �]�r $��q�V?�sd�����G?T[dy���d6#��n�disg@�������kb�)���n�G5E�ynJ3���,V?�AM�k�v���q�t/�6�u͞Ab���tҫX�3D{]�1�N�`�L���們]�r �r�b�0��+�y���ץ\3��dRN�H�����'�}@'��Yq�����g!�-��Lg6P���@��e��x�k����x�k9C:����zگ�A''��3�8�v��!��x:��r�h� ��K���^�M�	1m;zO��dPx�7jx�l`�c�'����ζ1�"��$�]�� �4������Q!�Ρ�v$�4����H��Ό2ރ�,U���lYm*uS�#��B���Pp�!����G&A�ȥ�z0����������b�-V��yA'0��'Sl��;�|.U���H,W�w�/���Ҭ�ɕ�˶�c�?[�b�;��y��mk?m��n���PK   ��*Z�i�B�� �� /   images/8f10cd51-b334-43ee-ae1f-f1b63d43b44b.pngLzeT�M���0�,��-<8���ww���	���!@��}yw�۳ϟ���9U]U�V���(��A�  �ee$U �,  z���r�4'� Pd%���������͹�	(I��W\�k��gk�������������X��{F�3|y�D^OW��rM��˻2���)��X��s�)>���JD}��͹��c�O-����Y�ͻ�n������u�IS�؃��������1p	c��@kh��x�m@V|���_M���Β��� ��Bt=6�O����=�� �lWr�>�x����>f���;����rb�È�)�F
��~�'?ke���%��X��_���r++q��/���9!���k&��d9��^���a�ӥG}d�'�)rs��d�'nϼ@���~;m��A��eT��e���'>a9V7ם��ɗˡYnf�}���.�XT��}�t�RW�;<dw��� /�m������gl�1)�A�.M����ndf/��{��z�j���Y�A��G����03���<%�@9�&�Y :�h�J��ʓ�0�DhVҧ� �����VG����d�h���������4N�>��9���ҡ��P�,Z�曘����ÿ���nG����=gmsN��i��vA�C�7Y�^��N�Xt��'r��/�H�f�O�^�k�c���p�I�zl�U.R �� ����&hN߫���ZM[[�b̩1��[D�$	����7�Hu������r�dV-LbV>�^"Mo�Y��hvK	Ƹ�_���|�v��o��{d?��6?��ڽ��|.�#]Y:DM&WZT�f��-���)��Uiª�r3��)�����&M5��!�=�y�rUr`��5���qiPPh�v�˦ů�O��'.O��8�@qb6mg����<���}��!�c��<@�L^������ @����@P*S�Iu~���K9��vx��M椋�=����ڏ���Vd���R�t�X��2�����rۅ�R��^9��z]	�p;n�~ u͘��|�iN:�٘�����d?�����.�n��t�"ǿ��/Bpi��D_~Bn-�$��ց�v�Q���I�5���VrU�}	�[�����FT�s�N��;Q�bHy'q�>�Կ�xz�������?����t�x����ΰ�u�6��Bf����0r�ws��'�<�*Q�R��9_���H����8����{���f�c~��4�I�$=�c��4
N���;Y��ĽmP$����9�<0�E��<�{#���I�;¸�bL��)���s�QT������ a�
��@���(׫���;��Z5>uE`�gM4m��h���A�|�=��@C��w�ҞS�`���0����L��6t�)<���GM�0x�Q�e�g�g�_�g�X�����I^�+��9�B:.�e�}��^�&��D���+���#����9��z-�@"p_��8nZS�!�-d%��>-Z �������TDB���<^:�G>Z���#�K�8�Q)�9���5	@�Q���bw���:Q�>_�/�iڋ�� ���5�����@��.$ p��bd�	�6a�e�	� +-s�gp+aT���	����FV-��ly>�q�uیM�0�3�+�a����r&S2���*;	֨��r�+��b�t�����Bax���7E��f7�3��A��2V�$k�5��t7Z/W	S�];�Ep��ڑh�Vb���z5>����{s~ou>��@�z�U>�s�&x��)C7԰B��5hR����3U(��G$�xS���?�	�t���N�Yg��z��)�h��SAx���^
{ek�]��~c����W�b��cs���{n�e�S�bK��i��t.��v��g���QE��c���4X���;���6*_�Vܧ��kڟ:����q��lkKK@�8���e����r�櫛Df��E���`Ɔ���J߯��/ ��y!�p2��h�1VaY#Č�<�YA�K!����t���O+��s0��A�¢���I�����]P������a6�1θ;���]&���I`�a���c�(it19��7�^emw����^��G-�c):::^�NMDZ���Pu�;j|�Nh��Ǹ���TH��۸_����A�Sz��EU׽^�GCJy|>� f1>���V9/�fx��eU0���1� �Y��Pm\��s)MS5�8��pc��~���{����v�7�x�����G�Yh�꣏� yz}��ߵ�E����*��?<w�>t�?�R=��}-���Ԝǧ�q�R��8�����6�s!ا4���dW����L9 ����RC�.??�}��t���6-�����D�H�n��O�r���Llu����d.�jw�o�z�[o:���B���ۮ[�;q}O�a�4;����e�c�R��0�71h,'��ƖU잣ހټb0ٴ�M�KC����ͅ�.�wsDO:�D��|6u��@r8QG��;sʳ'/�n�y�>ϕ�>��09o���ڟ8��8r���KNݼI���./bc#P������b^��.�1uk��:��/�<��>b�c���t�JS�g9q�����a�Ց��Z�_�E�1q�i߽�;�(��}�8�e8�{�KY
&~������G���ͳ�r�i�l��Z���I�o�z�ȟ_w��ѮN���>�َ�#���Z�6�����ž�U��<ߎ��U�SޓGEO�����B��$N6S�4\�5��G2�R500�o�p�%��;���ސ'�8��Y�w��������V��Z^�����A��dy՗��4�Ҥ�8 !$��J�>�)�[풋�6`����u���s��@%яٻ��.�-s~��r5�h�9�M՜s�܎�/:���Y��6��OG�x�*��:.u�V�c��m�q�R��e02wq�~ m �޵ߕ���<.������������?�r#��άB��t��+g����=�L�?�.]����3~������x���r��چ�"���T͗��Jǧ*��»7�4ܷ'��-���}�p�<6������{��� 63�B?�4�;|�̿�3>��m;��>�;�������V_]��>�]��E����&���������jl8��钗Z����@����"�#�����fO6(^�legw��@�Ly�0�	�[J�c?u;n"?���S�����ڟ���T�0K���Y@��>y6��=�k��	�}�~7N#S�H�qǦ�~�2�G���]J�f��'��Y�0�Z�=y���d6������o`ο��ה0��� �y݁<�w��4�ho���w.����­痂<.q�F̜VS<�7ۃi���{�=Z�/Ǣ_����ig ��[F-�M�`k��?3���d�Ά����. ���[/9�>^�{\�Ko���������v��!��I.ڴ�5BE}m�����1ߠ�}��2��z���c ,%��%�o����N�/.�x�� �AEٞ��ogd�kb�?z���9��NRR����ٮ#W2xH�S�3�݉G���<��T�K��*���s�0A��kzG��yY�?r�����D��;9~~:n�XkS>gy����!��!�5�aS�%��AG�G�HL?m���~�3�J��'ǹ-k���z�i�km)��&��#O�c����:��	{8���Fw��B~g�������J?�l��ra�0!^�4}pLn�~Z%��R�jWx7�K��]u����S&������~����ұ�����I��)�Z.t^��R�0��6[�ys�������a�`�%���K�x�}�V�U<�Cu���1�Sj�A,�
׻{)��9?Iw%z����g}��X�[&^O�:�⾇Q�T�._�N�N����"���n�+�{��i ��{b��ڝ�x���i-f��(y+��������'��\��&�Fjt���P�ۊY���?7�жїy�rqq!#�ɨw�z�������oN��u�d���S�E<�"1�@�,��8�R�����>&��C�ZZ�n����n�=����j���O�N"��z�u��%b ���d��_iDA���w��[�_%�0��)�IC��뮠�Ye��^�C
d,U��r����9��ڲY޹]�=N��:�Vx����lrpUj�'�&l���(���b��1��~�v�/��lҷG~dQn�_��B�W�Lf�]zs!Z���(q9�v����=�=�����f
����b+�nT�N�*FX�$G�8������<k�������鱱�g�	�����;q�O�^�����Ƒ:ԩ'������µ�i��??G냄Xw
��e&�M���~B��v��*m�i��a���<�����p�9x}�w=�}xjm�\l���m��ϊ�(�4>$�����_��Y������L>�R 4Z٥o)C^ūV҄�''���-_��C�׺^|u�~�]�@�h�����Z��O1hM؄^��w�w���j �y������ �������T���.u�yO������j�-z����Cte��b������야��ʟF���}��(�_>K�T��|�NL�π"%����D�w�&��v�Od
����Ы?j;d���4�p{:l����^6��pi����֏^9�Ҿ�/-X�z�=m �M ȶ)lň�_���J����q��;��$��f?j5��Ya-��3�^���i<��刄�G�T��&e�_+�}W.K�@�����11�� i+at����'�>O���G2�"�/4�?=k\�X�[��N�[^Zp��Ku�8�M�eT?Ȼ��E��.J�ZB���5���;��H$� ����?��?��pW^�aT�hck1��yc�2��rE����v_;ۊ-k=
���V��c��Ф��TI�4�-�X���T��-�H��I\Qe��AHBd#����7td�k~$����Ꮞ9�Ф�l�I!��7���6iL>��1�;�.�w<��~��j�s)���<��7��q2yQ}���O�����uޮ
oh����m���]������#�#��E�p��n4�G��(ҵ�"��4�l��?�_�Qa�ח�Q�H�457���;v'r�*.�Z�b��'�7hyeہ�C�o�NZ��
ګ��K��z����vE�>t-q�5Y~��pt�E�]b��?�RCP+��[4���o%�4a����{<g�V�OhU�V��^���ڤ'n���AT'��RA
��	Q��(5���4a�;��k+�0Ub�%n�d�}�����Ԭ�I��>-E$M�K��`�*�nu7�F�iY%D��i��{��oy��ll{:rg�ںqQ3�ߨYS��[d��X)�6Uz���m��i̥a�'�b�U�©���ǿJ1Y��i�W���8S����Ї��7fo�����F���u�tHb~4[t��W��N�u��!w&���J!88�(^kC2�"�L�] f��W���$收�����,���9�:�T� (3_�
�&���<ϫ���aâ�=)�����)AK��1�j�=�Ø��n�[�<fr��;>����=t��8!bO���0�Hv*����]f��e�_=��`-��`��9��jK��s���zty��h���}�ː�]����jT��.�T�.v�\m����?�����ɎK�*�W}�f��5��v4֨`W��~�irc�I�<��Ԑ�ET�'�I�Y\,����S�9��$Us�Y'��������6L�
�z�
�>�r@�`���,WW�U�:��z�*yx�� �2�O�B��	��ydy8%x�~�Wxh�{�f�>|��F:y��Z�zp҉T�<�b���\�0��B�򈅁lzKcV��A��T������-������ߛ���Z� m�<,��/�B17k;��<��`��yw��p����@jDfwC�#�W#��������_=��+0����'�DyҜ��O���#'�;�&,#�~%L�ef�[ӡ(b��~ �{+ʯI��J� ~9��9%[�����?lk3�Ŵo�+�O�n8��ޯѤ�睹����|a�t��CF�u)��t��ܤd0��;W!�X����W53�h�+��n-���-�V0��9 8�m��0�^R�%U.��i۬)�՚26�4�����K�ִM��y��=��av	�I���e��h*vxeB}��i��*R�O� �RF)����2Yݸ���:@�UӑRd�o9�*������4B����ꤿ*���$M9��-,4��ӣ��1�Ru��A j�0�������!��:�)��-u��p4����/�i�y\��L]�� E�;�:�IP�6�畔��vh���ޞ-��"YR�9�p,r�h�\�����* �m��⹩Fՠd�lb�%�{1P���0V��s3�p�T'�fqC72Nй�?4���
)e���6�)C�㶉�o�5�(,�"r�7i(��Zj��u^]5v2����iQ$Y�L]Е˳�5L�����i�}�!� P��v������&z347��&����|{��췎�EH�J��!���x��,i7�Y�D�r`F��f�HX�=`���R�|�d�r_�o����i�&�<��~?�(�4�R(��![*QNb�5h��7�.�t�g��2���ڹ�Nf�E�g�`F�/;YmVda �q��)mB0{�L|��=���70?`ͼ�����ڗO�҂?�vo���Ctt���� �E�_ɯ���)17p&D�nN
0R�2��wߛZ��=���`�*������d�����Ďk��n���C�6��"��A:�ȁ�D�԰��������T�Z�q������}��U�E���1ӝ���ֹ�me/L�ߞcD�HG�Y�)�D��ݏ����#��<[wsg��P;�9�bV�5�fF"B�(4�tW'�wԇ��3S�?�7�'U&�T��X�fXlO�gѰuT螃I�k�0�|5X���6E
`'�p/��8Zi��1�CǝR����::zO�WH#UL�B
 x��ԉ�ԡ棟����Lŧe���hfX��Z��"�F*"�@v����z�a>y.W�I�(����˹�P��h�(��'!y��hn����o����ݛS�����s���ۡ��)��k����H�����߆[���d�n��e��W�N噈)%`Wx]B�;R�=�g%>iM���zt�����f����De7%�֋~�A!}o�gbejk/����4�X��^��h5̢0Ï5/'`�����"�ZUn�xoܐU����lW�c��Z���Q�*��qe٥o�5،p�<�P�n������DRhQFx�������\]�9�9YW&�W�y]�;`�������B��v�:� �O�aÐ3��/5�O���~c
�痲�X�s}�%��β������=ƃjq-���^{����I��,�6+��.3�H�����z�]�}�|=PZs����i��c����D/�6~��F�.�tWyb��j������{U���W�fIY��2PC�e�d�V���a��q6 _0�'��u%���P�1��|�9�4��Q6�����	Z���|��K1��N��W�o�)Q�P�����2�/���!c|,}یTB�ڙB�@b�W��ಲX]�;I��!��K{�q�b��g��%�
W6������j,TV.���ѽ��Sҧ�w�$��G&[�h�"$1�ՑtS�ҥ@��D� ��sm��'��I9߷�{�?m��Vj��PF����i��m��}�������bq�Uq���ӿp$%{@�I���H- ��)�1����	x@@	��܋ڢ+����n�����B��2��IwH�i��9:�G���\�v�8S*��(5��\1�|Ce�H|���7G-M%;���_����*F,�1�����Y��Z�ƌ� }:�]�E8��z��ɉ6z��C���L9���8�ʶ����}}���F!���^�9'��k�Ӛ��w���gO���������ؤ�L���I���� }�6�u��Vi�`���pqks��u=�I�/`M����9'��ű��/�]g���,r��T�r�}��J�{,�vK��R�����tPy{��\�p�%���\������0p9�Zd�C��3k�P��v_�<S��?����V����}]8q�i��;
�~7�&�� 1�F�3f��K�q�U�i��1�p&$�w��;��^���4#vkA,����
���A�0�$�+�^�����i˗N
��[��������|�1�jۨ�~!�*�ady�x�����:(�h����.=���9Lё�-)�^h�DE�)C�+1%͟�\�)m%܃���h��+mF�F_j���֣���f/��<y�zy5(�_�y��ƛC���e���CH�B$!)a�8>���a�}��N������eH�~4��.n�b���oSr�
W�I4FEgTa��>�38�/cj����
����s�&ec�/k��x<��Zfs+�a��mc�h\P�ĠHt�S����]�����h��1I�w��Dl��A1WH.Ф�ͪ�6�in tg�n4lm�2��U�g��>�e=�pL+1�8&_�6�x*ޗT.�7yl6���ymb�,�rJ;u�b�~6(Zfok������C��S���dL�?�0�PIǯ�Hy�/_z�' i',��q+���bG�R�M�@��SŖ�����R-a��w:w�֌���Tp�C]ع��c	p��r=B�wy﶑>]8(\��%Wb�#z�=��o��w�2��1�@uD9"������@ �z�L7�=���:��*�}�H�Q3p��#
:5|��ǌ�o}�4!��1�2�&Y�aIǅ$(㵦u�����WA��NFbF��F��ޟIy��(3S���YC�oM�8,(�����FѼjL���<OY���
�9�BKV�gEAQ|?�M��Jj����O�n�&X��ϳ}�t����0��;��C��#�V#j�O�oh;��7HasR8��'4��*l�������iB���$���C��\��w�~f��`������?S,}:�> �����N6��d�-����[6������7���
v�3&)��_>�<�{����f� !��y:�5�=����OƃJM��W�Y�u��=��X��b4}���9�����%ܪ/�ŬE˚A�n�̀��vGD�L���PV����A�Ү׻0�v��;䄿�#�z�U� �?Ĕ��\���m��b�7\��Wh7��b7��ock���YG��Y�2��]f]9MB��=��R�p'�-Gq�Je��EoϏ}�|h��w�BB)-�d�$�|ˏ�?���
�k��b�/�ֿv~�IF)$��Ć��R&��.�W���T0ĭ�[B�4�a ���S(RH����7(�9��$q(a���2����1�.�~����<�:<�����}��ڣ���jQ!��5Q���Ќ�Ah���*Xq.s���� ��}��=��5�0�@l�?t���3|�G6���-��I�}�èWqcH���^�C�wp��� h1�:vF��ri���:A��#5]�I���?��z���C��I���|$]�b*�E�ᷣ=�q*�|�J�;8)}��������`���r����� AV'@�CQv�, A�f�ڨ6g�M�!ruT{�e��<��H&�HG��	{�i��[�Qd\�\2��-�(���F&�ޛܦ���w��F.D��~��,-�-sA��:؝���g�D1F��g2>�� +�޶�o����}������|%C�9D���q�77�*��f�1E֠<�N�+������\����'e�2	�RΓ9�$~m<�����Z��q�l����D}}L@�OG0�\��αHw�̲5�yRPZ%a����Z���^�J�� UP���B	������3W�[$����f%Һ35`h�Y�׉�> D 1"N~�H��S(M�1���S�szx���Y}��呠� ���ea!m��[��bNV�{"p�g� �N����3o]>_��U�R򝲼a
�u���Qxٗ�\�՟�:�$ �g=��;IԨ3�_�����C[v�!��T�H�N��G}�3��1ք������<GF���~,5q��{�J���4j#�{��<-"��?2.F�[MZv\Z�+� �m|v NæD"ة�� �=Ϫ/�p ^~��Ƴc�6�fO��5m����L�$=�@ԥ%:����\�.6�Z
��YT��|緲S���˵�|�\�Z8�_���"�@��dQ*9�3��U���?ׯQ��j�c[�:�R��VJ/�j�V����<�)�1o1�-J�(ԀɡSi�7��LF쇴�S;~$�f�Kncr}���Z��O���ɐ]
N�v���8���j�'�5�ͩ��~d30vn�U�z����T[A�M@�dS�L�U�g�26�B-����^�]���k��W�q�d�5&eJD�;�7pB�C����#G�5a$�#�-�+=M�Y�X��N���#���x��	�͇ۘ��`h�-B��9�F��n$ ������$�j�����]�犗F6{�����z�ŋ��;�o3�Q�Q"]�+)��tY�$i�u�eM����'6���hq�oq����AM�K F�1�`xW
��9�:�
)n+��t�j�2��|ڡ%�_ݍQ�Ԉ~�u���F�{�"ҔC���'�5\���C���OT�TVh���R��t�������`�4n�A�Ƭ��F���(���E��F���ͽ�r���-y�������Q�U�g9LҰ�(tM\���*���]9��ttO+��L�L#��q�1�?/9bbH��ܢ���<�O��8h��H�[��P��+��
$����O޻'|��D5b���-Umt8vO���X��q6U�x��<F�A��E��訢6aAἹ��~��q�6fZ1�ޅ�Wd�����ko�@�p}B�V�%лQ#��$J�.~ʎl�_k�22�5�4p���9AUB	ʐ*�T@]8Ux�����<l�����~w1�DX5�\�Fb\��"�oyԺjٔ� ��6-��r������c��l���l��۞J]��+rҔ��x�F�I�&��n��x�Z���d|�@�Jې^ORO��M�9"�i2��*I��M+is.��T�l?z&����!���=�9J��o��ג�i~%�w� AO/� ��btiY��:K�h�����c�z������?A� �Zv F�%�U+ƫ��Az�SP�6M9�^Y���H���������N0P<�b*���Ċ.��_�N��4*�@� M���%A3����z��k9�;�ٮ�����A
Jie3xX�G��~��딂UTH�P���a���)�8�B��{�Y^Y(i����p�m36�p%lY�����Ȼ�x۰� �� 2DbyYH~���k��7��&��d��T�r��M��5��s��f�)����g2�,�����܁x�.R�FǪw�RR���5Md�m �d~WM/R���T��QW�c����o��'�f�*ǖ�g���o>S�q�������:���TBJ��fBV�Ck�}�P�u!���GP�"(�e�KK[�\�2��-��7���]	��p9;c(��k�x0-kWe��PϚ�ŴH�O�;���w�4�������^S!w�2�"ہDX�r�j�Y��y�l����P���`����Z�ȥ�&;���¤��SlM=a{En����Z��8�ڈ���sAD�l�^���	�LV�PϚ��&���B�A�ߞ#��C"��į'H�~m�#�ȕ6$�ad;=���"�o��|MX����:]���+�s��Km|>��V!�KpeU�d↏�G�+�����3�6s���w�t_:�h|�k�#�����
%��@�!��X�i�t�|h)KB��"l*��m#� �wL�����o����z���nOs☘sM�ټ��J�% ��fڱO���:K �r�� �`l��Ih�v_�.���x\M|����a��-L�hnD���4��b-?�]�Ҥz�����w��^��Mw�� |}��ӆH,�*>�T�f��W��	i5�g�d����U=�zܜ��c�h�o���K�4~tm�C'> �'%���v驠����m/bju�Pn�~_��v�YB*�A��=�%�<e���a����]���!�F+����)�i�"�G���MV��g,"����_���W8���ॅ��{����V��}>�^��{�N��y������^M⍦4��\��q�e�������Di�A���7�:�)��D"�*!e�R�2^���[?��곍��a�����B�J�鐆�B�U��3o��!7ۄ���Bo����(�2u3����f�YcH�qv�j^�?~� �\�g��H����B�$�XiC�䷢��aV����<�Q���z9j�8珳��Y�����wxC뽑I���ٝ6�	"��z}��.s<�(qj��6����0�ҘS�N�EY�F$�V'�|�	4AsO *��)��t	��O��,���� �F�� h�|�w��D�;0�r>Ǔ�ߩbU�^��ͻ�(n���n�B��{�Vb+\�B��L��b�Me7� �;q�Sˆo�kྦྷ����W��l�\H>�qir>ƻ��%zߣ�����1 ǂtRF�9V_�-ԳG%2F�S!�,�\$Ǥ����������L v; D�O��������t�c$(��U5���ݰFd^w0�Y�k�C+SJ���||�Hr7��ݱ��$��8;���v�~���gg��wuR�4��0Fv�Q�to�\ 4��Bs'�/i���a�������s�aHt^�C>�R��@EE���j���_"�A�ݚ������>9;9U�%K�ko�B��i��!�ZB��G^�lS1��-g�?W�|��wG`���hR�Rw]!t5RB��
:W���uӯ׶��W2:a�����-���"�v�6�R�* +�ڔ�R�P����j��׫�%���'n$I���%��Ӫ!�D��>�f�޵����@�r���(��qk8��@�����V����+7F{�" vw�'B� Sr��~�5��gh)��-�|eA	aS5��N*d0�����9okICz�[ku��[�ɯ�7�UZf�@@)QR���4v��u��	w�V�A��B�8<��]*�^��p���?Ev�v��1�fcf����G�R� lF�5$Ɖ�����c�R=u]�Lo��X���w��n����̢��I5.{���6����:����}��V{�u��C���� ��ry;��o�ӭC���� حw�R1I��A��-ؓ�4L�E�!pU�ݰ��-����P�nz��D>���}�L�S�����!�I�̄�/���&�1���ܶ�I������Y'1`��:�����/e0Q��L��V�� c�l��W�A(S�}��'|��P�Kkg�)9�D
�#VǠ�SV��oe�tѦz������G)��ՓY%e�ӸU3��~�^Yi������X�?F��9�֤�>/Jͯ�C{�r��?��^b��l;�`���}&�Rʿ������h�ã!�'BS�]3�Ѷ��" �7`��]+��H��	&쌺U:n����q��_�z{�,S��ވ'���L���5�>D���m��s���SM  �HZ����զ��}��o�0�Jr.oyL�r��로�i��ù��'@F��G]^������Q��z���Z���+�R�^,����|Ao�;�75!���S�qR��Y������<d�]����c!_:�Ƙ�b���8ɼ��o���$޹�Xf�|I/q�D�6֕��?�H�ُ��F<�!��?Ku�2"��C��=�q�t(`<����J4��l߼��jR
�B;<�[��4$�ˠC�ȼd������W���-�Q|���>�{���~���)	�j}�q���O�k���U\D<�UĿx��+��;�����Z���$o���']�9�^G�� �]^�0�S����rA�35 �5�n�.����������@=�uPE��>9���ǟ ��C�?b�B����E2*ɜ�;""�h?|ǯ����|�c�럤1� 4���_�1���3��v�l���B��|�A&i#t�0��E��tQ�4��lԊ�����L�����	�Y�dHet�mR���Y��s�*<l!k�.�}S��mұ��s�	���/�������fR��� �6f�����+�/�A���޴��-u>2�E�ֽ��ƍ̆R��s��ٓ`y
1S�}\(|��?TR���X�9��'G��"G2=��/�U��/雭V���h�G;b�h�����	tE�2��@)��?ñ�>�1ݎ���_�!w:s�����'�s�\LIf�l��>϶'�=�\��\��+���w�����h�1�����L��axga p��}����B#�UQ=	�|���F��	<\���B����;����d�w���[	��\�b"]t�;�toD\��R�.�ٍ#�cyT�⊼�,b*�\dK0�@M�D��j�t��.Eqxr�\�b��?��u�����%��R!�L��(�ْ��S�_�{�� L��ԁ ˥x�~�
]cx��l��/3��`,�/���Lk���7Hl�r�`���7Z���D�T��'R�H扤-�'x�rac�"��ą�2w	�`8���5JC��W�Ǐ�Xq�[�'�z�����>+6�M�	�Hń�lҟ3��~}<c�2�U=��W�s3H�p�9�EnZ}��hUM�.��uSX�7p�mW��*��_��D�2�r2b���h�aW���ڊ��0�L%������^9��Y��ͤ���E%���2���f��A)���A$����S�`;%O��bv��s�M���p���\�A7+�5����=�����@�{�`D�N��{�C��A��*�yD�/T����/�_'��3LThRL���X�?���?pt��K�s��L��� �[�b���Jh� ��-�U&�{��L��
<�9��x�Yҍ恳ڀ5��#~��Y]VP��g����5�0
�i�,���P��Sܨ��_0DdN
��6۶����8>fe�`�Z/0vUz`n+�׫\2��O�P����Zĵ�x���x�b�b�#p|�����?T��
�eP8��7�˷��B�c�s��>�틢��lv��#���99*Dn��c���5c������]��Em�Af�\Y_f�5��K5�;��?0��3>�����@��.ˤ����M�[�+]{������ߒo(?)a�t�Mq�ܚ'e��y	���$:�����Ԉ�?���%�ϮG,Hwn	���_��U� 6Yr6h�W�u��_�FH�|�x`m@�[���p
���w�yf؛K����5@ꦘ��� ��5�I]�;M���_ˣm։R`��Q��󸦘��g��IDI�w�ط�2ϜZ!c]��@b۪0{Y��?w8�Qt.U8�l�W�h�B�i>+3t���̯&dM�<��1n�� �B;�������3Էkw2_j�r.���U�0���U_�ʛ�Qj|Y���H�2�g� �D��R~��z�oe�*su������dw�.6	��w�k���B&!��Ko�����W��U���t�B�eC����:$��o�ҙ�9�}j>8EhA��|��^�v|�&nQ����AF��H���%(��Mk�L����_/�h�����k)�9�kz�1Q�Y>�W�7 ��	�VLU��!iؔ�Q��
X�/���J���<������d�t
����Z�mc��"�1�,Cx�:U��=ɣ�4���Ri�����#��P{<������+;�+�"�$Nh����4�#-b�#Y�N�4�X@�]�W��gh��.caf��������	��i,6�~�\wFF��.��}G@�2@b7 �P�k�.W�\QӇ�g��gJ��J�	2v�ŷxT�R���?oJ\�U�#Z��O�^�v�L>�l�����1���h�H�kcժ��8�I~���,��T��	�а/�>3�nQ�qx�kO|��ƈI�;0�׸���X�_���d��QJ�?W̋g��)e��sR�Ý`y���=���ZXUA|1^^8��h�'.�Ǐ�.��F@������3�*�H�, V+Qv&H8���2
*��O] ��}��#?>^��4�����f���X��%`3��b<��ր�)H_���a��ϐ����	tÁU]�h�}�1�}�<d�~	V �f��W̟&󧢚<)�8�H��������d��(
9���������cl� ���%��Ɋy���R��'v��nVj��e]m
`�p�o�=*G{�O���́|T1v�{�m:��e����TiH�4S��x%S��ȯG��Gb7!���� �hC�B��kAb3��f*]�$,5�[�B.?��X�΁��2�'�$�� ��NX7�|Q��QW�WZ�����:��x,�C�uD���%�BW��t�k���e�b���8T��^!��;�R�ߧƲ�_߹N� W7�C�'������Wd�,�ި��D��	;�h�j�> �c4������bZK�(*0���ɛ]9����Rl@�	���EL���I�?�а�?�^2�t����n�r�T����}�"�`�<����c,Y�j�����J~�)��Q�'�E3��AV6HTpɂh���6�мuC+o �_s6J˒ݜ@��C Y9�@��C9���ɒ��L�����1;S�L&�� ee�\���t��E����  ��1G�*�y`UO���TX|?r��������|!���CH�M�2��%�X�f��g]��IVc$]0�0R��N�jA,�m
�gP�%Y��N͝4���O�9�w>ר��غ��8�yN�b�8�e;�r�f���P�k�qw O�L�6Qt�a
:�m���g�n�S�
V�m���nC`� �^[�i�(և��Z�i(F�o�B�7��#X�E`��>�J36K`��,֋W�T�X���M�q�1F^��|�T��/ +���E�#��Y3�&M)�5��J�⺁��~'k�������ՠ����(@`���,�P�5c�3X�� ȩ(�RB��9L:���i#_U�d�A�c�	�κN�\`~:5i�O* _l�N��(e+�Ya"���5Y_.��ΐ����>9(Ͻ�G�J��a�+���~8fD�
���ܖ�:3^x���}�F�X'X)����b
S��/^\-Yx�N�q\�$�MaNk+���jq<�zT�.B�+!5ç@�S�0�Rfb��t�Td������g�kqj�ͲV/�7�`A}�}D�Q�U��-���2���5_�B�3F�c%���$
R�Pˇk���Z�4,�U���@3;��9�R���-	�pL��Mcs��:�e|>w=#�*jM���ǋp�U��v������H�?X)��p�è��bi.<sl��y�>����#p�Xo�bj�r{�*ɉJ7� #]�9>�ƈK^f�(�;^A���0k�2�OB��r&�vQ��*[��H�WU xT�饦���+�O_����!�v��,�ۅ�(9�>|r@�}�t��*F!
�W�FS7��8���G�k��+MO��_T��o�v�پ|'�k��zɾ.`uZ�P`� ,cA
6�.d�?l�R�3�W
�'<���տ,���#�������B��b�,=��
�2��V�d$����y�Z�V�Z��@�+�2�ݥBQ��z��C7��}����(��҂�Xe��m�K��n!�^��eT`U���ѫ����Uژ���[��2G��qP~a+�㶩�T��^�*!�HY�N�q�{ J`�w�p���5�6k,��}-˚��
b�\V���֌�挲��V�ۘ5h)/��ZYh�hP��_�oqdW�g�Z'�R7��S�5q<(�X��׍4�C'3���r��� +�N�R�|ݏ-�!;_TX�z����`Md��_|�Ee�r��'&Y��n�:u����Wy��-J:Q����)�_�˒��d�,4�TtZ� M7�B�e���yJ�B,[?����
�͙5A9���i��c�	b��T�FRM�-s�\��:�"�z*8�;M&��\�\�<����F���[F�������Z��s �X/ZlX�7HKY�+�*w)Hze^��b�<��Vٴ�b�(-�r_�F��2�}:�E��b�X�y��r��5p#�����ͬ>s��ȇ��Lq`@K`T@%S�TW0���0+��x&Sb�bյMV�S���"��6��N^�]j�C#�jI���t��ڮ�>�(�Oo=���G�Dmه㨲�p�����.�Ћ�q����V�XIJ���L�⃸T_�l�Z����w+!��:����ݷ_/k��E]]�;A�;��XX�%E=u�X���暱�vS(@ t�t���l��G:P;=,,.b:^�դ����
n�ր��XI��
3N�)���ِ/8{J=*�hz,#Ş#��%ކ(����3֋W���VF�?Vdǜ���		�Ե͔���c�};����D�%��7*�,̠��X��G �$!���y�:�uc������&�$+�ZIS�~�
̸�Z��)@;�4f����m�s+?Y�Z�L󩹶	����9�M�5�j��]c��X.��c$!�x�<͙%k�U��n���x�V�8
�߁�Yyj�������2g8������V�eh��kz�L�uZ*������/^4�`Z����rXi���Ƶ�^k�3�+.�פ+G�i�>8���$�N�[��_!����k�/Ӗ  �p}���
�:����\v�������֙ҏ����gd��nd��-C讵*�K��/���\��̒�$��[��V�k�`Zl��
;׭\(�u���;��z�L�!F�:�nB`���˙��b����Ђ2e�!�_}S��D��G_�!��nSF.)�)���5��+6Y��4X�pG�����#���w_�Nn[�"=hL�������(�C�rg�T�S\ӳ��`���*e�<� I�x%�	��4)�W��G X!�k?�	�@ -@NP��V}���<HTX���+��-֧�8��hV`k�a�HG�ܗ��2�j���B0ՆE ���s{�bE",6�Nahi	X���ݹn�,��`�F��W�^��!(���^g*���^�JZʲ)4�B�U���gd߉Am��ٕ�s��#"���hLJtpE�/5V��KV6:/�RqM,��~<��PNCa��o�RV�l@���J@�A#G���|т�h����	H��5PF<SM�,�������I7�#�P����\��\T��J`b�%�=˘]�X	��
B �w]w�`�s��[ڜs/WKW	M�O��Dr��'-I��V�4�������f�̮�NJU�~."�`?�c@�Aַ�#���TR`���T0L�Y�j_�8l��ޭ��8`}r�Q�XsI����J`E8�1\l����-l+�����b�X���5}N*�u���j����%����K1���d�3zч�!!���#�0Y�w�p�,�Ղ6Oi��6 ]
k.N��ʂ������I" �<6�Z��L�n���s�-�
�0�̻uj�q<��Pc8ll�qC�g���mކ�]7�E�8XwyX�h8����Tj9������Mā��gԊ�I"����lG����J�������X-M��s���h�T�iu�mZ�݆m㔈AV$���2r��b��m�r���t�<�3�<�i�~b��A��b�Rl�>A��҆��gÁ�5��>��Ql�^=_�~�,)W �IksS�jhD۸W�6�4XO������Wn�j�l������9m����m�k���\����k�����$ �� ǎ
�۰u���f3p%/��l=IW/+k��u�Ay��7�H\�� ��:X�u(�r�Z�H�`p����-�t'd�:�}5Y��jFV����CP�Uװehv�^��UY�)ɥ�V��A��J������,QU`�Xc�+ �$� �� ���Oi�2
U�p�4�7O�2Sy��.<8�g�VǕk�ŏ�婮`tZ�+��S��k!٢�C|��`� �@��~�}5��s3��Rŋ�,��P�]u�.|+,~��&X
䞱f���g��XAH';�wd�Q�3
����cj�,�DQ�w^�FMk@mP,"�!c<����e�:��X��k=�.�����4�\$=Ť�x���X����F� sk]�B���Jv	�N@��%5H0��;+W��߼l��s�:���D�Qj���C���>Đ��6���Z"Zs��%#�f��>�E���FA��eI�&�ߐ��_q
.<�c9�\���8��y���Ե�1�TA��*i�C����3�z��k�)��a M��`TK΂�%��H� V>��1+�4n-����9뼢0&��ӭ?�%%�,_$k�S�8��	�wA� ��x��9���A$8��4�b���e�#�g�Vp�t���ݼ����QR�.T��s���rC�Ƙ�y��^Y�`�� ZKB�KRE��甛y,�Sg���_���������۴/j^S�v������8�����^V����k$�-�A���VJ)W�s�j�V�~��՝�L�1���a�44������<|T��NH�D�D{�$��d *ۅ껁+���\�Ǽoi���6i^0W�Η��m�C����/�n�Q6��}���$^a�H92�4�X�lI�b�)��~������y\�q(��*�˯�h�]5V,�G��b��1Vv���g���dV^
�u,�X�9q2���H�CH���&V�.�I����?66`Ąw�,@۱V6Gn�R���ɪ=�&�K�#X�qX��u�R�����<�"J��b��\�j���Y�S�F�x�.\�iX��ŀ�@( Q(Q�=�[0]��&I ����eTg��Fq$ k����{E�,�5
�v�(�h�<���ҁj51t�`�su�kR�	CV(SW��h1�Y(�=��T0P����"�P���r�4&3Ha��*4!XR���f T�Xs���ǚ������:������do� �C�D�%�ë*X�Dh���A��JENmr��i���2oV�V��|�ѧ�?�?)�d��Q��}�ʍkW�k�^�L�+1
T�D(���±=��~/>2#Y�<S����x97�ɱC�e!r���k��ű.�AR�gU$i +�OM����ٲ�l�FPK��qS��k�VɌ��j�"��D%�Z����z��RF�_��`�%b�0X�7�s��#���ʯ��Q9/!'p����)�c�$q@��/ͨrԂ�����d_����^1��Ɓ2�A>� ��T�d��%2c�rI-Y ا+�B' �b�@9hn���L.i<��<_g�+dX�a�fX��+��X�ϱ���V�*�4��H����-U,���#��B`��u>^���T����U�u��d&;�����z>	.��+��J�����5�pj������2f��X�A�蹎 ���O�&z2�m;sb7M�7</��і������6��Q�(|��Ȃ���:�JP����`q�\�.�)��v�4jq�B�9���P*N XA���ql+Ś���
��<��&9I�`O`5�bZ �RB�] XP��'@s�{B���UХ������oEo�zTm��hi���W�El��J�9}�d#p�W��c-��'��<���8rR"Pz
��=��0�w,2_���
�f)ۯ䥙m�2��UVâo��"���ѧ��>x#X\�c�߃������ ��B�k��:�ۛ�j��Zl�5�h�r��)B!�8zH�,Y"�g�3��y̿2ݪX�Y�~�{@��u@�>!��hr�K�\����r�a����������\�:�Z����\����m�?rT��qi�OK�~��>�<k�7.)�
:mJ#BR.)�P�p �V�o��^���BC`�N�n�4�X�n�"葃6u$;a��kE�UK5��cx��
A�%	���c?���Vp��Y"c�w��kP��ᜡ���r��>�!�h����I����������L��@px��Wɒi��^�X�G�J��1����U�=��I\�M���Z�����M��[�y�-�A��}ʍ��]�-"����P`Q	����+��-kWI=I\heX�(c��2��� � �t|�V7����m���!lPe3d���R���0�L%�j�q�~�Xd��$H$����9��
rݕ˥�����Ɖt_Ĉ�b�+;� [�+����T<�&u3������w��]�N�-�����>y��y7#]�	<WZ�$��>�;���"sg�D���������O��^�.���[�b��\�|��b���+|���
��@��UD�ۡ�e1�����Xw�te�"J��]'��/w0�r�+(�Z�֛5�U�p-.J���,VsP�zZ�4��Ni��nd�����7�m ���L��H���TZ��Ȝ������8���v��sPt���f�C�`Q��=�	���o���F��B��� ����CVg�����	�8&�	p�<N�5�s���o�	VO�1[E���8Y��EbYy,åqB��V5:u#���m �Y�?�DՕ�3�d:\:)�k��1V�fl�1����@�mj����gO<#;���x��@�)�֦�m�|�Jc>���7˸,���`=N�Kh>:SO�I�~�$�v��U�*L�g�G# �n��� U)��K��Er�j���U��ɬ@c�x�@���Gv��w���)��Ye��56D�6������p�MUkW����$İ��C������:܃PV�>EP��@��މF����y��FBz:��d_�D�P�D����n�e�R���Y�V��f�-�
� >�	p���KhXı�}Q{b�*�Xd{��E˖˴9���M��K[�*�` �P�H��"v`��7���s��g2AS����g���X���5��p	�pIBbu6���moȡ�_��X�-]����+S �S0gS����p��*�N�w^7�0���T�W!�!���ҐD$��|��c��L��Z�w�m��X/}�6Y��LAL���g��k�Y�k����!�^j�p��k�f-ل�H-4�dTp�DYT�m�h�j�$��ѩ1�zɄ#�.�u�b� � �j��Y���XM�k�'Pj��#_}}���A�h���k��54��\F\�,>�K�Bq:�$o�HY7E�3;� e��r*��-Zv�`�}R� cY�2��ةV|!�A�A��#-����_�� ���k|O�A����Zt��1�(&��t�D{vX� V�Ka@����>Uhpm8f���pQ���{���Z������N�
5t�k�Z�t��zH�W���>��"�+������.�m�]�u�p`��Fh��u�s��<T>�!�JE����y�v��!KV��ًVɣϽ,O��CbM���8>HC�ߪ�1��,;V<�u�.R��{�X���6ut����<���g�k���W����o@��?+3�}��(C����EmWGД��[*�l�'�rW�,�>,"�څ��{-z�;d��7���
 �2�c=l- ����[sf-r��m�k�NO}軟��]���C��M�
�
)L�`��N0�����k�m��hy�� ��j�J�l��?X$M��A\-�RIZY��\Slvsaw��ZM�<�B�pS�#J1�(Z�Z%K��c���Q���!��h�;MV�L��A�$"�l�h��T�K�pu�Zi2�wC*J&�t��d���!�N1�\�=!-C�%�d"�F��IXX
,0�S�Vn9xtW�\��W�ۊ/�j�5J���n6�X	�ȏ�3�K둬w�L�.&��p�)m�����Ú.3ǐuZd����^r�A<��Rr��8K+�����Ș�q^e�Xˈ;�1'2���}83@L��~�^yb�[6>��;$/�QP&��\�f���O�2/�cGTC::/5�(����
��؍��    IDATV��/�&/��$�钫�>���|��Jf.�¼C_��Z{vV�w,�%����ĚDU�:x��Nv��矓TG�,�����j:�5�<	\���hU�ү^bP-��@�
�NX�[z�B�<�#��0�]�`�f��˒��%�E� ��L�ILF��ylO�"���� �q�<�R��Y��x-V�y��Ȑ�k��:XG�H��A��P9)�ϭ��Y�\1�^IMc�[d��̝0�����d�x�L��xp�|V#�.J��X�G˕��5\�4�s�K2X��@��`�&��BP.�їN�K:���c\�3�-�.eX����B,�{h�R�Pc�������I�rWV��\S=���������j�,FUx8Nt�2�c� ������n����$L��9-�A�S\X΍��iar�1�����z0��uR�iFV��x��K�^��%h�d��W� �
�,��;��^�v�<���˒��Y��Z�g5�8&���Y=�p�SF�����=Qz��`����WHӬ����7�m�t����AG59v�������~{;Fp�/D��X+ -�#=2�ޯHR}m��rh�&Y�
O)�s�Ni�熜���{�%�"��i]=6w���ַ�?3f P��G�TPPSxKg���>[v��q|�Z���}Q�����)FO�O&�� �J�B���
�����?�퇎���\�~���:>�U{�r�a��.>k
D�X$Mp{F�='��
	d��Dg�V(!�`�|
έ�$($˗�U�ucU_�Z`���>}����T{�sV�\���,(Q��!���aѕ�+�qPwG�OO0�ź	P>��*Ȫ���<�y��2��k�V���P��B�ǩ��#�8�Q>���Q��r ��A� *zD�>>eƈ�����UXX�܄��>4�A�p:�5r��܅ b	�l߀��vB i�4>}�{@�ZV�2�� V�C0�&�<��׳���b���ˢ��"%ٿ�,��:u�* �vyr�.�4�k�C�S�}hh8�֔���{V�iƜ-P�}�MEaX��](��j��!I�6���PY��C񘮎��ʋ�J�@F����I����F �vʢ�K��M�)�[s�u��6���fv��c{���´6�Tq酇�p}J��]�x�:ه!T���Sr��_�]ģC`=�����d,V��Y�c��Gs�f�k7���Vh�K�ȴ��|��z�D�ዴ��G�Mc*�L�z��L����=P�w��x�,��.8E�h�Ǘ����3�ފd��4�!ֻ�Y��/���� o��U���_2���@PΙ``
��p��hZ:�R*-�K`��hq&�u���� ��O��X܆�H^-��ل����\���J��*M����|��X��Z�O�{��X�ly�
�����m<����t�)|;�
������Ҙ�si߁��p���p���n@�BA�	K�iq�o5$p�바N�� +}7�B*�1X��vn�[^��0uf��h��Ƞf���.X��VS�Y"h�������I�%�`�Bc)!� ��7e��J띷�! tJ,�6�&h���ձ~����G��?0b�����-ʭ��z�c<��Xyj������)�z�*��e�bh!;I�Uٯ�VV�$��h��rF±s0~�_~��x�;7���9�u�-�(`��Xs�X�Sd UT�J2r�Xc�ƕ�`��`w�� �#�5c����h�e$�3/8
pe�4R�(�P�
�H�
4(,1n��r���jgb�lٱ���*�G`��p� �R �fo�&Pu�X1�}�2�Ӂ�Rv�>yྻ����֙��9���!���ɞ�)(�"���y�</���e��+�e�Jyĥ'�D�&�n�8W�����6�m��8��ԿB'�#h�+�^x^���#�0��]�2��:��h���Ħ�)t5�W���V���G����Qf@��#�A�H=
c�'G�]b�Z�s�{�DC��"|U"���\�V3"P_qމ`�6�JWp��f��@�VNR���@�������f��X���� �c�J��Vj�\�ͫ�e܃���(���>'X}�)[E��&�w������h'��0Ӓ���C�@7�<,����4ku��k ��
-�G�`�i��>��0���92�p�wmk�&�kݘ�x�!�Qҭw< �ʰf7�xJ�Q�SAÊ3����"+;��ti����=#+�fm���l�V�0�j��	Y��m��ڋRs�X�����̚91V#-������K��&{��H#���Ʈ�3�ֶ�2����G�WJ+\����]�ڲ9.(��њ��.y��j�~�	�X	�0o�#�������1�*�t�}]�.� D�L� ��þRYV.��{��؜��(�ܗU/�SE3�n	$�&j�z?L+u�BY�+�(]m��%inZ�	s�)c8���p�9�����}���K��B��	�q�i�Z��y���Q�Rwc���5���ʅȨ�i�>�a�NZx�p�ߝ����@4^�Հ��n��Ms�z�6?v��܇��h	(9|^L��[�,�X���B��9�tY_WK��k>G��m�^�m��w\�C���:�$R�9L��u�бdz��~�Zi�L���ԉ$�G_�$��P���=`A�+�<���[�J�E˻0W���ʀO��N��&wM�V�	l�A���X;��V-��[6JX�y�l�j�\��r)�f���p�;f���Kd�
Z����k���T5;��������䥱�Xu���\@s�
� <L�B棈E{ڀ��G�9+�a��aI2^��"){���������=�5��,96�ь���?���,�`�e鞊�yT�Y�Q-VzgjY��	)ixF�5��x'X�$��5u�q���z��k��p׀��`�=��b��~ZcNA���C�ç�x��t�d;�
&8�_\Zid�Ś�����ϒ���u�F ��V-k����Ø%K�B՘�4v�՗���&�3'Yɀ�����\�M�A�����P��f�*��G�Z�3S�{�yه�y�o�^���b�8�%���dAW=���
\#f��WL,6e/�)v����G�Pm����+��i����,Z���+V���,��g�ָ+�F�f�4z���7Ui�\	����ic���Ȃ���:����k�^�x5�	�Np�Zʔ���@^���!d!��^}�Y4�'����s�Gڐr3�k��`j���0Si���H	�θ�RObI��Vr��+��KO�=���~�jϽ�^9�JLi��2Kz2�+�&�).ּ#�ቨ|&`m���h!~k!^��΁�ri\�piH�T>�SsY���Q|q��6r]	��ZdPz��.��}Ҁ*8!+x�`�lyF7!���
Ej��bmBY�)t��N"ۣ�yɥa� ��&�N�6le�U6 0�(c[9W��Sc�V�9�Z�� k�^Ӭ�~뗞�n
y��"��	��p��L�]�ӈ%j<��5��q��;��gй�ca�Gt�3�>��?X'�_���J2��a�(r�b�~�r�y?��g��OH�C_̨�ǆdJ�۔xE&7E*�Á��)j�|�\��"l�����s�1,OJs�Q#�����g�\�y&�U�9� �@�`�$�ʔmɖw���I��c��g�gw��>3#�e��x<�	��lɊ�Ŝs ��Ρ�+W��~�9U�
���$ ���ltwխ{�=�_x��ق�:�P0���
�G��K��� %;	`]�:Vn� a�<
�K7e'�N������1U�V�� (`�`]�k���Wv�o}���̸2c����G^�0�����*��Q��=C����()[3�h�ᓲ�8̱V��8o����Z��v|�	3R����g����c�I��쨎���O�*C��:_��T��K�\)�l�K��|� :}dȱ���l�q��>G���jX���
d�y�jR����u���Z��Fd�Һ�u�[c�ۢ�Oli&z˄�ޑm��v�-���M6����Y\��Bc��Z>���!�+5�B�>K�zX�X�k��������ڭh/���F
����Z��_-��P:kC�Ŵ��l[G#:�0���d�|n�v�Ӗ���(������^��C(��q�+�b�ܞ��`��B�V�h:�.���+��85o��a�]��j���2�
9Cz�dk��s /X� �B �jM�l�/`~��m�\6_�R u�Ճ"�l�VF(� �K�X��
�N}�e�m ��u��#P�/����p> �24��6�gf��H��wnG���S�m��ĨL��K�O�Mݫ/J��k�!N`]�E���@%�2�k�!�&C����VO��@k�5��
�P;x�Ӗ}�S�}õr��,�SӘ�$�?pFkb`�k�<�w:`��|F����������X��<Z�(f?�m۬kͩ��g�q.Ka^�;g`eh��97M0���X��ˢ=Z^+X�Tc�?uu��+T�����iCK�K�+�&R�^U�����Sn|r D��b�� {e4c�/����B�x��2�r�*j�f�����@K[���������-�Ju&U=��3J��B!Bnx4N�F��<g�+���!�vŊ~��-;%�vU0��}r"[�<��@��jj�~nB��ٵ@:YC�$��X������,pG�K�v�X"��[ϯHaM$1|:����0r�Vn��O��Eٵ�2y덗%�%��m�jy�mô��%;����d�Q�5]���8�&PB`�P�^�E�V��G�
~��C�;�
��>WO�2��f����
�cU0/���c=��b>Xaj��RC��Z���B�QD�8'b���R�K"'��R�t���b�.� z���7���¬G�#;X�*��	�_��A�);���JsR��2�^�"�ߍe�p���P-(/Y.��3Sv�9
C��.8XR�
hg,j����� �C�`�����q�y�H�֝�,4��|+K�6��6��cm��C��=j97[RV�e����X �5�k��Jz+Vl����;A�C+;�y��f���>Q_�Q����ֆu��ɲn��r���	�gi���k&J`en�ީy��Y��r~��]K���R���6T�B҅G�A�̛�Ǟ�\�T�e�0�us�b��Y	����h�0�T���ܺ�2ٸ�S��:�����G���`O)֩C��u&�r���4��q��;���:z��B���Xg�A�`�����+$ùq�g_��\�m�^y);���ܼ���M�L�����.��4�f�U�yM�B*�yi�e�˂���
�-��uH*iz�fp�
����u|���
��5u�.W̅3+�hPZ3U���.9��{��s/�Z�ׅ��90(�(�递�2T�
��/"Đb��kL}�ׁk=�H�/�T�hA��!���6Tn�FV���5YD����-�������;n�������$�R��,�]T���jV2���+���w�u��P}&�9�Fu�B�m`��C�+�������k4O��*�X<�����t8��Yњ���N��
����B����/Տ<��q�Lԧ���\�z�`�B b�
��f$�87����d�2dαRQ ��X�P��鴀)`��U� �X袖��U�Dè(8�R��
�����]�>�v[Շ&�x]`y�f'�؜`Y��8��hEk3j-�y&%ֿ��~ +��B�.]�q��el���X� ����/�О��B���W^���#�����~����@ap��\�bh����T�=�k��e �5��ֶ5����q�' ���l���Ͳ�3wH��WN�=b�`p={�	�Ql͛K�p�����*���s��ҜC�v9A`M��ԏpp<; �Ax��F�h���h��B�VlrO��5��J��z/�f�n&�
�A ?���;�4>�1N�n� i��5,{ r�{�/z�N8Bs������!Pj>A���=�*�sa줌�'��(ڿ1:��ru���5jg.��(�]�2MV=��<s�]а�4��!��a]*C��N%�i!���U$�p�&�a?�R��~X羈�r��X	RYл`z`�@��B��^M��h��<9,݃hWD?b�F�{��!��zu���k8���@� K-�2:U��p:-0HG�0�����|Z◯�}ж�Y���JO�?*��+��'ق��s���{�X�kV�q (Ix�$/�2���k�l9Z|�l9�%'�Oʐ��n-Wq��x7���}=^ �݇Y�W����9��3��j���-��p����}�<n��o�U���5̎.�E"�����8���v���uD!��C��E�tէWIk��)6���ŭ�[���a�
���&E�6R,{�7JI��-Z�{`��s@�
@���ͩ!nX���p�+�<vv�,�}�ۆ�-R�k﫯H��>�[�C��މ�����^���O�Lv��;�n�Ӏ�l���̜�X3���\*��y��V��c0t���-��	�z�HT�ԕ��T�$�2!�vm{��w���D��D l�̱�������r����4ު�}��gmA���ms���{mR�qr3��îOAJ��5i�C�XL��:yI��`�xh�3
&�Z	�l^7?��5�gщ1��9�"�;9 #ޒD9�=l-��)��M3�	��_�in�����P9�ީ���=(�R�,%��0�ݵz����6#�R�K���B�k��/�s9���$�Q�+���xL���<59"��|]�CC���S �ɂ$�K�UI7�,R��,�s�+��k��%*�OY{��'v���$bұ�r��f���r����j�q�j���CɅ\�ʮ77I��#Vn3T��ڡ�s���k�X#��F䥩��
F�k,�2�|B��F�a���yY��ar�}�N�z8��F�p��p��\O�
�[��=��u�����\IXYn3�B�>��L
�<#Y���Vp
����y�)%����*Oɂ���Q����*�U��с��%gmcmC�"4('YD�[�v��j6�����e��2�l8%����2��c%��}��QW͙��n묇n^�xq+s�Q�駠���݋���F�Mc�c�=R����eh��P��h2���\E�q��Mq�1d�E�m�	I����v���i����CE��,���s�f	�|�8�u�e��6Dg�˚p��h�~oHs�G�����D�۬�yY,�p�9��P� LJ�NX���B�'��FC�S2b9V�	�k�kU����n��L]]3�zv\��ژ��ו����Gzp�lc��_w���[<��K�c����m��8E���]�Lk�<G�`ͯ�ÅȄ�peN��U`�����4�kFV=b��tr�����e� �1�3I!�_Ǟ�'[�i��@��0>�`�Vn���C����j׆G[b��h�lGn~�wq��YSM�d%�G�HM��]r�� p߮4"- Г{�Jf���!�Q�z waM�7�ճZJ�{�����w���厤$/�E�V��5k$�t�����2]�����:c-yŭ32ك������еW^j������y�+�7���X	�}��$!���TaG=k�6�V.��3V�I-X��l<֍�y�ȣ9>&2�O��x���Vp0t�͟a�;������`S�����*jA�e�+��I]Qk� D<XS�C�8O	�.�*=���
Π��d5�R61' 1�j�%�ce�U�I�5��遵�{�"l�����Q��:j��&��z��i��#̓X��;Ģ�ę�`_�c��C���Vi��z�h�����Q�3ѩ���Ǻ�9�J�Zt�y��3���������0b��!11�m
�X1#�{�=���.�������3V6�>�3����æ}�/�1iB e)�:V+�aY{9��܆=V��4p>E�����    IDAT�K�`-P��H&=��A�+Ԛ���HetT*ã����
q�4{���G�锎%���}�D��@:	�ԛ��g]��10�V���K�t��Y-��,�2%U^�P����a�>L�!��H��Xg;�>���X]8��tg�YX�^M	=
�B��u� ��]���d��2����EYF
��d�m����9�I�"�Cߤ5ʒ <@ÿn�*��|+`a�Y��1 ɚ��&�r��X=r&�,�wzxl���?��~���"x�/�,\/�Qy�I���XQiZ��|���Zcj�O@��P/��1��"��
���c�"�L��}oH����L�Bew c"�;_ዄ�P�U�* ]@s�Tt�=��44Rjt0��{����%䈦Pnӿ�
��^"����&���"?����s��~���pI!�`�Ğ�
dV7�AL���B<�Y�D'��3] �r ��74S"4um$)�#��.:�
�y
+�ek��	A�ķ>��\e��>\sȺWO�$H|M�*��؏X?������ȍ�V�
*1���$C(�~�Ȱt,��}̉r��e��h �yQ�H�������<f�xT^r�C�+s���ĿZ�5��d�iXf�Pb�V���`8����UO�,��R&��
�{< {r����һ�*I��]m��l[���zx����;vO�>m� 	���T�Vp��k����HJ�cmV[h
�Ⓗ��Z3G�S7��exߛ��"T����\�E���	��ާwU 4�`3:��z�lMR���X�h(<��HXZ��
����X�]'�e�}<g�鷁u6�6ﹸ���o^NSg&�0�N��=Dʞp	�Č�"�[eԌejط�oE�r��~c�+%c�6��o-a�Ȅ�"1�ͦ�6�lqV��/T��#՜v#����r��ph�#�X��:KfFg�'�uZ�%LD/��c��+ü5� 5vvE� %�0ze.Ρ��.,\���^U�������}
�����-��@%�O�O�)�Q�\y�b��6�3#������uN~%�(.ѻ5�
������$�� �2��%�G=-�6Bĭ�JH�Q�8@���e={(��о���'�%�~+1�K�$>3�� ��,�$mp�FP�aI�i�Z�*��''���	���כÎ@5�Vx�\.酫] �׌�p�
�~6H �Ѽ�����6^���X� �2�P��y�6�b��j3�o\�:�x_�b��9����K�6���m�4R�B���J�c8)��fc*����E���
�XSV���4�zF��6����9����*D�����nB�hD��m�:.>��q�l� <��!W
�$.2��cS�ϴ ���\�I��ʰ*��A�S��s0�˖M�=j����y|IL�-��<��5`VmR�rs :�Z>����6H��r,V��KR��>!�.�\�
3�|%�#ht��@�^�u� ��������4�"�B�W��#��i03"�Tj�w;� �a?���!V���cQg��U��3�6�-�xZ��TGe�Js��Bx���0�i&�گ'�E$�I�DS��ٯB��K���P��B��֠v�[��g�.7�ͳ���c^�-wq+;��y���ztS�9W����B����"aR�2$���E"�wm�A>��S������S/�C��. ռfWJS'eq�^����}ɍ�c�����w%5�\��SIkL]$�n��m��#����j���j89��R��*<L���c���~��(<O�K�{�ySxL�փ�m� �+�9�BJ '�	O��"о��w�)��m|�\Ds.&;�~�l�F�{<j�S�BQ����������(ű	���D��+E k>�X��� ���ܛ�m���Ve�+ul\U�1�Z�Ӯcdd���H����jfy�OȦ5K��k�#$�	�?��+r<���(>�%�e��] +[�i)ƣL	�~	5��/Y(7mE� ��")y��W���T��O���H<���k�X�}�<��D��h�lFm��sqk�2�+�KA󐚼<����-V��~b�W!|�NiL!�w�
T)��w}�}޵���ͽ��@.U���$&�BrH�K
]9����|�X��:�b�g�'`�Tuc癪ۤ�����ؼ�+��X#�i�c�fa���D@- �4ɺh����|	�a�ٺ.grF��pѨP����
�R�`��8��Qf+��(����H�U	���YFCp��q\��8�z�*1������k^^�K���		i>7�dl|/?G���mt�P~�i�00�d�s�S�p'eբ�\��R�tI�v̡��+��g�;��:��u����.��l,���.��"r˶�r�r�'~.�����(��9&#��)���do*�S7c�C�Y�)%��:��x~�pq�%���R>z��땑�'�U�*��(	�x��$��4�c�+A�X�7y6��\B
6�����v]�T#d�o����hF
��z쵂r���
>+���n����7:�%65��q4�f�*���(��F��F綑��)7�����6Ϋ5���p�z���
������R˯�H8y?�T�akOF�xo���R�H�*�J X�ᑲ|"��p��)~O�}D���	�t�Y�|�z�%P߫@j��K$9���Cr��I��HNBr��,�|6]��kW��nh!N�g���Y(4l;啃�N�X�
9D���7�A��1/R	Y�r�,Zاy�*���zu1�G''e�aԏ�g%/��0+s�qg��q�%0h�nd=Q���S���"��z����k=d��O��|v��(0g}7�~��-��W��%��!UQ�Hw�8Zf��C/ȡ,��hF]T6" P�j��G?��ÖU=�����nx�a���c-!���^�w#7�p%<����|�&�<nc	s(�a��6:�Dc��8#�mPr�;�G���۠m��c]l!8�0��z�N��˦����QGC�=K_S�������d�囤m�c��q�_l��1�!������3f"�:C(��s�V�a��*�@��{h���5�zq���H[X�zlD��<��OFl����"@EܟV�g�g�䆑#��Ux�È��17�qM�h\Ƙ�ge#;`���|��a��1���|8��!|TF+(���+;�Wg���k��'UV���X�c=`�a��F��U��tx{�}Ő��@Q8`��j��]Al�X��~�1n욼n䐼vO���7�4����)
A�7��vՎ�S?���/�*�z��8I�yOU䝣�9]�E�b� 	Ӝ������vE��Ƽ)����r>n��T�	��C�����҅�e����P��ٺAv]��(fr��y8(M���<������o� �7�ܞ[�>7^̢mRV/_ ����҃s��B�l'��	�s��<��s2V�H7B��΅Z��(�!��U�ݻn�I.�l5» �BQZ���A�$j�x�9rbRJ��z:��P+C��`gz���D�Bn��r�f {�3-^���>o�I\��/�ңǼ��o�5�r�[�j��xE<�)���{M�cc�Z�y&�*�i�hA�9O�B��.�Wo�NR�ce�B�P)��>��>1,54B���� �t�գ8?r��C㚴Vc�9�	L2[��"�3�F�!�}'���?{��x�Vy��%;>"+W,�<�ri�3v5�1�5t����'�b�|	�1\M�zVx�,);r���ذQ��(�������P���
*����(���c�}!3rB� Ԟ�H��;��Rv��}�Na:?d�2]C��F�w��m V�pc֪�2�ڀJeD^�l�����a�����}��u�Jf
�V�P��6�2�W�çlh�<P�0Mu�6�R���ƞw������Q�*�U!������:�۬\�1�g���h%|�L=V�\^��s X��y�+Co
�x�9��:�"i���}�4�_�F�dI� 
��IH�ѹ��B'�ڡ,�0`�+u="C��z��$Pn�����:'�G��t�gX��v���6��*)�Iꀕ�_��8�6��f�=�Yu�"�	[�qQ:$Kz�w� �â!�H2�2�*2	���>�ٽ�Е5���x� ;.[%����FW.�0A^3�D;)����_#6�Ój�����䢩ʚ��l�t�CC�tAJT� KS(?��5Ll�^��,�B\> ��yt�B��GX}���Y2y�\�)_�m�yl�jq�Y����W`	��.ݧa_ߓ���s�Z�{v,��n�.�LX�{���ɧ��B��P`�A�(�>��E�Iq\�R�l�@Hcǩ`#͎�DmaF��}�.�y�F����T��+W� �ƃ�Y������O��B�L�o@��@��̽$��+��(+/���&y���奷�"���M}��q@i|6��6D��FO��.�b���r�՛e��pRI4l0tu�ަu	����I���jڌذN�Wy���;h�s�?�a�K���-^;��t,R��8�"��V�uEi�������v�����ȴd�2ȍ%���}��
�-"JX���o� �u�2�sAÒ{��\�����o�?`m�X9!*[�o�I����V����* ;����+�;R��h�:��c�-+�ga��9�uk�>��_T��]�w���ln	��Gd [�w����N�� ���#S �{�� @E�u��L����X#*n�,'�8N������~�Λ��))�.S�`���E9\��l��@���=''�'O�"xlqCb���dוеxR*�	�.� B��┒���Y5�#c���䱗�c����K�䋷^/}�j���ey���'s���o(2�TCȡ>����{��pp�%.!�����UR����,�/�z�+\m�gL�0�?x�%92�0x�O�b��!�*3�[�5.����?}��@Ъ����1��G��ǥ� �27Uc��Y�h.|��g��\�SCw�!�<&�c���o}�+r�����W^����=.yX�{��N�@?������߭  U�e�6�1F�Q W	k���ټUzWl���: �?���(� �s�iWNg�6�/�s���3��0��z�6ٵ�
l5Y�Y��@X�!d�۶y���\ ���e�SEzD�V騰�9�+�q$!Y��������b��S#dQ��KX���n@�z��~�u�tD�ٶFA�c�@�RRǆ&�D�&� F�[D�T�E��޳����t�ݥ9y]�����Gs�u˱�	さV�y���f%��G�*.|6`=�	�Ѽ�o�>'Ұ�������i�*\��>��`�7��3����G�%�PpNC��"x�c��� k�yS~6=V#��O���;�2	^P�5}���
&a/&�W�A6,�D��v&M��u�T8���I.��U�������W%�EEY�������mвE��Z�=S���txz6�pH��"�:VNʏI�d%	��ڞ�|���Ѕé	8lTh��2Ðs���el�%��"Ʌ������H��*�h��'�A�BMk�¢�$,���@�b��/��l�hHF,�!Q
ϙTk:E
A�0Y�8-w���>�ʔ5�}�������A
׀�7Z�cc�9Q$��[���γ:�0�gcj|�� � B�߸���ҵ2px��IC	��7*l��R����@������vF�q��ƒ�lVA��(��,Y�A�.����+���$z� |Iţ�>�z��T�5�2�3�ZȠ���[x��#%p�U�ǾQ>�^�ne���;��Q�� 0�S!/CN®�I�K`	���Xn�Pg�XiOf�ӈa�����V�ϙM6�FUU&�D���q���p0 � �(o㝽� f�	�Z&DS����:�@���h��3����Հђ�f=s���7%+�&�f/�*�T�p�c�5܁P�6����c.�mg�m����6ru>D�?Y���ȸ�T���\x���2!>�����I�b�LE�K$�blXw違cUV�!��J.`��"��鳜��#��0月��~�\�9Թ��ze�°l"�j�e�*<�Hz����_?�":��{��\������6�rk V�&J2=M.v�Q�R-�K`Ȏ�S�'^ h�n������]7HC����9X|()!;1�uz��� F�>��y��}"h�qn����Ҋ5<�4Ƶ?�g�R��R=x��HK�����ƙ�<9��DR���M�%����u���;��"�w0����xU����ųd�u��O#k_ShƞY
�.=�_������*ج*�(B!2����u�4�TKZg��|��3Z ~�ZtH�r��4���HV:�5��z؏���<���\��:��Ư�P�,��AR�e3*���Eg�n���Đ,��uWn�=�4rlx 2c�Eu�_��8"��>����W��/׶sgz��cU���n]�Zv�]�b�핔�2��T� ��U�s]���=G��[	\�"�搶��c���4��$�c���ֽ3\��G��$�;�G�:V����ȱ"�p�n�C�of��!qn�꜀�Q�ˁ3��zT�::����~N�Y� /�{�1�7�4_��X5�O�AH ��Lc%A X�:/s�۟�0�9l�QX���EY�VC��"$��p�'�Iז�H�=2�{Ht-�w���w�xa��q��^{��ܰJل��RE�%=M����Xp�z�Hg����ß?뀵"�-��W�@(a�
B�a�j��J: P����N�����}o�V�)���f�L[�QB7�M"��-�29�x�A�3��5�0�!3Q�<��~H�@�����OqASt��
rS,E`>��Bʵq8�5
���,w?7`e��*�`n|T��A
{��{���c�,x(�u�U<������/�Y����*��C�|�
��1j8؈7�����q�o(�RA�(�yPD���^{_���(Է0O�c�����i��h���.A�D�+: ؓ5��H���s��%��x�N>�JV��~.��T���7ޗ��{]�%�b�5$�i\��z&�U=z����"w_}9Ȁ�zN���u����(�Hb#~=�[��3���4"0\C ��)X����s���k�<l��Ȁ�&��}���8ZS�m#L��؇��<tT���T�a�bb����y�Z8�ǧ!1(���U��0t���-Bwy.S֪�h�U�b�
><���ʞ%AǺ��F?�,0�����S��+Cq�u!��T�%�qFA*��z�7�<c�Z�q�m�,?���ѡ�E"��Q���}C
�nL\P�?�e��|�Z	#�J����(7fZ���"FaѱjR���g����5�tQD��Z�)`�O!��b@\�b	��I86�<�H�_G(�w� XA��U97�j�3�\i4�������eBؠC("TN�9�
��Z��{�f�e͕�-	@��{ y�cFKc6��F�<��V#�0��߬��<Vz��<tA�<���v�"Yԋ\v�ќk����]�Q�0�Ql�.8>���P�2���2iG'<�H,)��� �n�3rm�
�$�� ��֟�q�#�ag"�(�2�X��[�j�e,vd��sEY��~�kT����l�y�Wv���e�P	��:�Ӳ�e}�+��V2�<VF�j�q��*wm[#屓ҁ�=��rXs��Z[|��������o�~C����SM֒%2���eYGkU)�r�3�E3�FXn��#?���qX�x(��aql��p��Q���j�-�6{έ�Z��E�u4a�D=9�؊)ʠu����wx@�K�k+�0\��ԀH�
�K��c���!&����I���0Y:�4��7�  �'Q�
�ËY���H���0EPs�X,���^�1 \����m��͗���G��vz]\0q�i4Y¤L�_�$���O}N�L`S�b^� ,_�mX���    IDAT�,�]E����XJ�*b3�X7s�̷&`�����N��w��C��K0=��	����١�HU�X^Do��zJ@ e?&X�w�7�8�ٽ��8e$q/1�j�gތD(eR��j�*����� k�Ck
9���!��$�K Zz�IZ�G��ע~�oqN�����f�w.�'�~	�n
s�ĸ�ш3���
|�@��m��� 
�ٓ�Ȫ��k�i���3u@�
q�э<ourPV�D勷]#��z�ԍ��U�������i0^�}H���z�a0�D�o�.�kU������8G��x7mY#�\u��ƎA��Deh�ǁ#V"��Su�������S�˾A�j7*N�|�:�BEdln�Z��y����^6Q�<s(�ӿ�<p�,7̴�FC���q���CXYLO���P�D	t;�O���n�d�0��M|��+���Wo���� 	�drXgm��q�ٽv��co�`�nNx��#�ڷ�-���`-��>컃��)�Fz�k�GI.�?����Nklh��NY�`��� `̿t�u��V\i���'# ����im�:��Z����#�!�HC�"��n[!�l]�B�j�2�	$������X~��������`�������w X���Re��b��5�Jd"	a�H�O��ݘCȏ��9O�_�n7�����Z`8�a\W�@PtLI�i�Ϝ�,��ԣ2�o�p|�����X��X��\�uZ]��H'G���Bm3�+��5F ���q�g���3�縊>�o���f��i}����z�8�R��W�0$ɮ- �����(����t@�8��g��Z�f��$Yd���I�21 �&�+��VE]���[��o݇k����#/�ok�g)�#TP��7�}�v�s��;�r� <ް������B�?�][Q����V͓����?\����zS>D�
�i/�Д���I-!���	��#p �	�ha�"�x%'ف#R:�!�"6zJӱYV�r�}rL�@�@��<;��k>n�1�t:���x�0x����2��������~���Ł�GOF�0��L:�ʰ_�"�X�x�2Uj��7���}8��%��=V�����z��`����z�|�r�Ԃ�D(3Df���
_O�}<�C ��#����8�s��	L�u�R(������ΰ~�,9��G�I5��\!�[�}
�zZ�f�{[��/�r���c�!�żj��J(n.��y�d�������{����I$!v��ĉ�}�g?� �Q�Ӄ�֠��FG���-_�a�o�{Q�����Z�s4�q�׹:����3��:9!E�S�����s���8�\ֻ9b�ץ8��>�qP��#n{��X�����&:�`�&���N�� 0��4ܘ�l4�Pr$��������Ġ\
N�n�J0�IO��r�`�=�������_~5�5/�ޠ3��FnF�}�5��D�haRnܴZ��&����̓p�HP�5���� D;���gO����zp��V�al�uP��5S��>��|y����ź�U�j3�;HuG1t5I��Ou���KGd�Ax�I3�۾MCN��YV6���ގ�\��<��o3~QX��q�����gu���`w��aaG�E�N
�5+�O�G-��J"�FoQxy9-T����sc!y����%s;�b�x$/1�J`ݸ��a<z�[�A�r��BV s-$Itˇ#9��?��Z�s@�	�b��5eצ�ؔG��I�Xb�)�=��`��������(>K��e	��S�KgyJ.nXYS ��[TrΩ" 	��)�P���������R�����c$��#��i<ޅ����-[�*���u��E<� �Ƞ�����3�-@�?���E���]�y�lO����sΘw�H6x�]��rkm ��g6fd���;	jظ&j���i�_�=oO��2��52K`���4��qa�ce��ϖ6!���_����xB�x7�5���2�p�̦�����|l�TR4��􈶅�z'�d�S8L��@u�K��ͫ%�e�����	3�`'-x��ű�uQ��z�y��c^�w�E�+��vj�ȳ���;ߺwm�������:���G(��|9Ӊ�z3L�Z�8&Y�I�J8��W�ʎ���߀�GE�ݾU7��՞�l�,��i�V78�1��z�e�/!���DΪ���LAO6BQ{L}� 2 �'.�`�l��j�B�{=�ȜE�M�ӕې!Ú��H$A�+I��`ڥ��XsC�����(�Ҁ,L'[Y����92Q��X�X,�c#��m�ʮ��B+a!����6�BE�6�� �?{��?��=*K:����"I +e�SU���)�Xُ��{/	V0��~���(�Y�1b�o#_=�O��gk�t>���<��YD?B�I��/�4�)�<���l7UM6ƈ0eʝZ��q�ŕ�g�bmܓ����:7��fe��L�C�R��cCG "�"�j�g���_���=$9��ᤄUswv{a+��OU��"�`eX��x�i��&�X��F�0ejB���9�sJ�7B`�?��nyꍽ �^��z�u�1?�%�߂=��� P�1S�6�+�#j ���5�|
҅�N85���?��/B%LY����a�����|��K%��!��"`X�`��f���8Ur*_�^D#Х<��k�Y;R�S	L(�:|.���D:�6y�h��{����0pc0`=8�k�J��:�^�;x�$k�P�+���������F.���x`5���"��ڨ���=IX���/�vX� n��!��a\ ��f�#s���C#Y��ϟQ����庭��v�R#�ع\ܚ�=��>��E�Qtl�α�$ju!{��/._��v�$��27e��r��N� �I��}�-y���
���k�F��:���7��x��������*���Ԗw�qj���	�k�#��9!Ц����$'s�͟Q�ћ9���L�h���iW�;c������+�kH |�0EB���^ش����'��[E���ڤ���%}�ٛ��%�H����J�1�^��}��Ĵ�c/�%O���rFX�V��';8����� +���ۯ�Rn��rD� `���(�9c���{G>W�T'��RH���O˾�1D���G�����R>��!/���6ICֱγ�zz`����ax@e��q��"�@����˱�_��]1ٱi�t�0Y��8���c��gY>����N?u3�3��u�P���~ k�+�FK�M�ؾ��5�I�;-�7�l��LyǈL��TaUj9��!ݑ)2� ��jY� XoݱM�_��%��G0I�"�-ʒ�h�b(��N9��x߳�I�j������n�-�k-'���նs��z&s��=�<��ɢ<Ծt܁'�~y�|j��e����c]	����S���B�u<���,
΋X�$
�/�.0�-�g�g����{&���K���w����vN;��7N����\�p�u�NØs����\l�N�����C�s�����
�d�z���j汒�g�M-�%̢Ս�ٍF�<j��P��	cm�a8/��k�]!:`�"��f5E,Xo��Y�N!�����+�~8`���:Q�-y�9���޴N��Y��{�0\q0�Y��D���ch)I�죹<B��ȇ'ѣ:�
��<G�#�׫���X�",�b +	P2��m��mb�(I�ƛ(�\�G�0U�HfP��!K;�r٪�h%�>�=,Y_g��P�}γk�9*�@�
[������9��
��ֽB�����E ��9I2�!k!I"�փ�z��kK�䖝p��D�	��
�`7!�P�5j�
�`��Hj����Z�%���h�����R���1.���܄*-_��E09Iz�M3���
�tUv)���!/�A�ξ#2R�M�7V��K�%��/����Q (sN�@ŉ�ł	r��rl��ha`���9?�yz��H�<!�5O�wޱ�˭6����GPA�����l�2�%h`��c����C��t�Y���^�J��GP����1\��QØs��'Y���:`��XcJ��W�<;C�(u�P�v�:��s.�}�NS�g� T# ű��wS�FW���G#��J�C��NN麯"K �M�=q��u�T�C^*����DU�3=V�k�:,�/�T[��΂32� ��+���ɫ;�3�mzb�sj/�=^˝�c=Q�ʑΰ��ms�rV�4WV����L����M�`<�"�k��#.,ɼޓǆ��[U�&����P�3%=дemwum+���3�,cI�嘟)��Z|�>I)�GJ|G?��{�s饈�w@oaXo�Л�N
0L�<�*�Xx��#��������hw=��LS��i|6B��
&)I�s�}�p��U�j�@c�Ŭ�$
@�Qya��Wǐ�MP3�4X�Ԛ��@���T�s��=�����	�`��B )K��T���%���J��2$ƨ%\c�*���5	K3���XT��$ �OK�<n�6��&����������A�U�L]y�B��5��&���c#�5��ok�ryڰ�k���5����:k����o�임.P��d�ía]�E:��T��T�B* �B�sR�j\��"#^˜>s��S���/	�\�Z2i��BaH�4��Y���v1�W�؃X�G��m2՛Tu1{ﹳ����fc�0HwJ����p�14�\���&ѸEZ�k�9j�m��X��y��}5�:+����s߱r��r$M��.sߥ (���}	 �/��3�wz<	��!�+I�'�B	Nl��L`��ɲH=L��km�� �M�����]����b����GN	@&�!���ȴU��<�����Z��/\{�N����f#h�����./Eɰ�����T��}>g3�ht�85�� �BN�J��hzǭϱ���KT�.Ġ�q���-0;����g��,T���n��zؽے2���4:ů9�l�˛N?��m ��^����G��_�?�t�����Mpϛ/���ϊ{�=�F��{w�y9����fDk�y��r�3pv�z"ƭ��jq�N׍3f���-�9K�5Ǻ R|����}u:Vp�]��7��XuI���W����9�b��o�D1AV����2^i��2b���F~sfؐNOJ����wM��Y�XQ�����-����]�ƌ~i��3�B@��>.��m7�ٻ(�����g�jF�3%�٘��D`�Jj��ٺ����/_��}ѿ@#�z��\�uf��9���sD�j��$/�X�`��Ǫ�y6��� �Ԑ$Ěӣ�wx��8�X,�l5�@� �8�b�LTP�wm3��-�z��>K��]����P�?����ZN��^~�����O]�ၚ%ܘ�zҍ�j�[��֜C31������K˸�~��7����萹P27զn?y=�p��s��p��R�Pý��1-�F~3�¤��rr.�ȋ�=+	�����)���
�+,4&Y����* ��b˾�-���Xg7���!n���v�����ׯ9.'�}\�#���3�X[a� ٘��50Δnն���$/�qo_{{Zk�i\�t��Ⅶ�\tIƹ���������C�荨tW�c�����-�%�T^=�dZ��������zvn+x��U���-��d
LNp����
��ąy4|Y베4%�cVz��\���;����Í���Om�j Z��,X���T:���<o
��o~�����W�1���= ό������;���is�
���M�X�3�5�������Ɲ�n��B(�Pw��JNb�k���Q��P�s��BKM�Ȱr#G��PV��T�y��s�N�l��m�`�Z[��q1���o��x��X=9Ó=,ja��>��S$�+����ib�,%��a�6�.��Ӿ湎�� ,4�ϳ��I�;G�y�g�����70��Oh X���6�V ����l���h�蘼�Uu�ΚWu���_��~���Qq�9X��Bz�Y�\�E:�6&P
���Z���Qm�Ç�U�}\�#� ֆG�Y����J*|iE�lg�mں>���7zl����i_�<�@k��?���u��;XE���?��_��c��Z�%B��ζ��U�@��>L1e��C �m�Q�-�::�J@*B����"�_�����p��u��w����Ӵ;5�l4��|y����g4�S�������]*4���:�T2����>.���<��u�X����k�*�֘n�6j�<�6o ����w��W���c�k���L��i���{��:���\�&�V�X)� |q x�lp�D��n�J#i<֞���Ha�e��e��K��Kd�~�����NAd}|rRFF'���r��A9|lHƲ��@O��G�St?�"�>�J��`�*Xx?_����2�[�K�X�4�ՠ8[�b���~��0���`҃����J#1,N׈s�������{��TE��ܬ7�X���X>^A���q�1<��G\�#��N�	$#��$�kr��t�Ev�)8:l��غ���}wZ�����'�+�{����J4��5:� * 9��0�����՘��HA�n\';wl�M�Ɋ%��IIW�ћ	|a��=��#�j|��d���r�Ġ���T+�/�te����wn��y%f���z����&�*r�z�s��Tw�>�LF����<	
@��d�2+L{8��u���?����K�Y�̘��4�O|�Z(S���F��gr��״G�j��q�Ã�_>�X�joV���k)�:粒 �g!1P��T�&Bl����T�ھ�(
�S���F���q�t�"�ʝ�ʖKWʚ��L�����G^�F׸#r���W�<����kʳϽ$���[2�Mu/��aY�-a/��i�*���"�ݛ��7�����~��n5LK�����\���9��kN�C��/�w�<S�ū�d�'�H�5K�膠�6�`W��2�́k��� U[��g���|���G��m��~�XG^�ӓ)�k�i'h�Gy�)�g�~�F g����m�{�O��W�>�Z�*'�0`� XSu`凥R�>6.�)���S�@��ڭ�Kw�(;6,�>�G��&��]6ICc�.�05�K���=��tt����cϽ,9(��Z�Z�>�ԃP`u����#�)���O�6�~d��1���&A��K:��/V[�?��f*���%W��<6�2i�������h����h���?��mL{.���Tbեd�7\>��^Ծ��A-� ��5W�>�hљ�x�z����N�b7*�:�[e�R)7%i4���' ���7�t�l[ׅn�g%�7E"���/��=N�"o�睜e_�Q�ߋ|=;�]�@���Sr�cOK�[�w��
�"��D���SU�q����3�XZS�A��ԫ�N<�B�f?���w�۬y ���Ͻ�ʵa5ޔ�L�ښ�^ ����(��25�>O˶�L���b˭Iڦ|9��4g��5�2���IzV�{��+9$�Z�s8u,}s,WyQ5j��W�E{T�����L�/��+���_��c5`M X
f^W�Z�8��(���܄\u�*��_��l[�/���j�����ͭzu-u�p�_���s��Y��f0+,hW���1�n�����}�=��j�~��^ڋ�y�>e�䣳�5HfOn�=Xc���әW���&��_���I����y�j�=�ImH6�`Y�(���~1Va�A�%G�H+?�9��xma�
6�]�YT���X�} �����Kc����6?���;4]TWA�;����=T��D���Z�QM�=��4�g�4��A�+�q^e~rXz���_��|��͒�E�P^�M@/�eN鈗A:�����j�(c�1b��NMh�MMp'q����Gr�������#�b���W�k��a@�u.S*��=[��f�,�Q��Z�Km
�-��ع<�㽾ل#E�У�Q��R}!��	� žΔ,]� �E����$<�    IDAT)�tH�i�T��p��Q��3~,3%c�Y9>0,'�Fex<#�\NA��n�j�&<�k=W�݅1��h�����M[�J ��
m "
U�P((ρk��"6�U�ۨe����<��{�X�ſ�;��i=��|��b7�P��A�-�j�m�������~���j=E��dOQ-�aȊlF�m�5���g�ظMe#�̤�ǲ����d��>���$�~v���_~O*qtjE�=��Le��i��V�� &@ٿ��:�-]@@���<}����f&��bk�X]=�kR�^��bMq�����kg�6Y?]O�s�j�W�#|��K�E�)��a]�r}���X��_6]�N6�]��"��Hk��P
���Az�<"�C�~���fc6Qg;]����ɞ}��	��'��V�a�C]��p�&?�i�[����F���G=G>�󛸈���NϹ9ʧ�s}� .�|��G O!�=4B�U� �UD��v ���%]�P�H'��c�8���S�'��d��e"�>�(�j�	��}�QJK��u]o���u8��\iA<�w}�[���@������?���9 +r��e/p+K�Q�AT�������˥oLU�����ExY7u���9Ғ�$έ*�P��&�bc������dU��?��r``RJh�]��Q�����l��<��2��@�����c�.@��r�����|?�p�n�`TK�9X1q2����k�
*8��e�?[75n���������� �̰Dc��7�f[��ʲn���~yL�l�U2��I�m;�i�����3TF�/}���`��,��QN����(#�,�L�����k���E����G�[����>\6��s@�a���PL�1�/��8�7�P0GO�
�^'�����ӯ�-O�I�s���йP�B���z�q��J�,އ�㆙��c���^�-�9��s>���;�Y�'ur�aU2X���ܦ#�{[i	6?��hM�M������=��Ǭǳ�S6�Q�+�s�k��O�%�p��q�XGX��:d+J>�n\/��/�^ k*׬#��+��'&�j��?2(o�;.�ܳ�����D���D�{ X�3i�/V��0�u%��0Q\�.����돾��i��	X���?~�x1J`��>�g�7\��ڥ}��u�f}� c��pO@��6�N/�~j��=�k������DtW�p� p�����ˣ/�#�X���$��`V�@x��wa�����	�և���KX1Ul.�b��c�i�䳓j0�|�	˦���ZtuhAˇX���w�1k�H�-cfL!�=��W�$�
�Ox�Ŧ��>��Q�{-�̍���V�:E+�ѵ�V3�(�,s���3��ـ���R���h�3�,,�����sty]'L�\�a��z͕���K%��GJ~�^YA,�p����<��J6�UC�u��� �m�|a�����#���Y$C٢<��[��/��	x�}Ka��2�R�3�C�H.;��p^b��sxo���m�a�|p``(Q�{���Z��s��IԲ����acFB�>j7�Q���N�ں1�(��OV]O
]t�L���H���tJ�SY���n���A�,k�/�k��&7��)�V$�����"���Y	������K�����g_�=�
�J��c�����P��XQ�^1�����/c-�X����Ǯo +@)!��._#����\�e���� ���C�@Ǫe��0�m���N��őO�O,�!�叞����G�R`UR==�O��9,XZ�de�5��l �EX�e��>��Sl8}P�Z�t���yY��[/Zh�J03����Z�~�ka�?_�gؘ�G� ��V�E����@>j,���LA�ȑհ�dk$����g����r
���s�q7$X['nXg�������3 aa|�XHV�Ӹ�Rz�e��u"�[�����˟�]�ۺIS'U�j�
��\�g����L&%�x���=P~q�H���������=���t�>��,��Q���Ert(#?~�1y��W$6}��O"�B^S
�|���\!0
��hA���rT���V)5FD4�����j�UY� �v*�\MS�{QI��m����*&��u6}���������D��4���@���%r�Xw����<��߭�l�[���jo]��Ы�½�{�FDq���P�O�f1q�xC��Cey���᧞�����{��kXG�9�j��,!+��ω3����ON��` �F:�h�2#�s�z����uY/�+��r��FC���9�e���!Ui�s�,#�8���3�} +=�
���ԅPm���6��pT �����J�%�� i.����C�nղ%���xHVT��f, p���.[�X��G��
�|7p0	�ƃ��oYh g�|.U�� ۩bMr �� �p�cmn	�
J�ЖO索�(�IC!up�~��#������|�
p�@8r��ڂ�*LH�<%�o�J���r��^ɍ�(�``uvv�5;::*�? G���qM#,��g__�~�x��<?������G����Fl,�)`&��Lv�ɳ��.?y�q96��P�!�N��s��ܨ���Kc�-�9?s��>�V� V�a�mx����&Q�����^�^�Lai����?��:�Pp+Od�1�R2w�6���s�g9���Y/��o�Z�w#�X�BjE�A����]��۶ɒN�.2j�� �kq>�k����&s�@�N�h����e��|)O���1�w��YJ� a*��5���id�n+c��[ �.N������_�6|����C������x(��\�i���?�U�X���4b�pqe{��}:H=��-"�1��.:�Uz�����ɏxB���7��V�G+�A�J�'��$ ��|4 l^EGL֭\,k�-����ZD�dvVF�expH�_۷m��Wo��]�|]��}3m6�ڰ&TG��(բ� �e��ɩ��#�18��LQ&k���R2�IC�U�B�X��ns��z9Gk��^ſ��灵U�ޏ�ϓ3����!_��gL�D���z����*!���w=H+L�&%���uN�;"�w������K�ʪ�+���C�7� ������L�c���͏s.�6����ݍ��U�w����!�����{tX���F9�-_�<U� #�G������nVK'ٽ0���;��0�����x� DP����|�h����ʄ�	��m�Z��B,c�w]&��x-E;@V�!b�����I���C7.�H�W>����[d)@?���b�&�I]M�bHټTe +{ށ�{=����Ἇ�x�m����/cy���c�5�ԫ'{���0t��n��)�X����U5xTQ������w��d�ʄ6�c`ֈGdRXZ�,��V3,ǡQ(��ӂn�����x^��Ag��[�fɣ��]V�Ҫq�33��Z���׮��+�H7��	X���J�����:۷1lp�UW�5;v�U���7N�z>TK+���b����q>�
ش���M��u`�(����ʘ< �xڄ�F	��|`��[(���lKxv?�2d�yM�+ ���r]����-�ꧮQ˙����*�T�(襖�����{���o��b�*Y�n�,Y�TC�EDR����y<_����M��kٚ�e]��)IlL �D'4��>904)����Jﲵ���L�����"����͙�]�P0=/l�X}e���$QI�Qֈ�^���kUi-��r��v�{���4���* !��o���먾G�	�ZB�KK1�#y�U�w���uհ�nr�҅���o�F��ջd9<Մ:y�F��`�CI\�ݻu?��l<�w��_s��$���:AZ�8�B2���?<+?|�)�
�Ra�(��B��(�œ�p����{�gfi_J~��w��
N+���NЛp!LO�Q�$,�/���iQ�(X��ט7jY����[G����U<܀�%��Aa>��D3K*y4W�7�k ��ދL6� ��2|��Lbcd-`�J!�4�ow^s�\��R*�<n�������@�glո�{k�b9�)j�9���h�$�F&��B���y����D�1|��a7��Βs��'ȅD�?�⻐��
�}�e��Tn�ԃ��� �PJ�����7��s�B*��gr��,] �M�O��?*�JU�K.�u�7JO_�^�P��X����t�u��5��s��x�$�2@?�]'j`��C$�x�<��a����TNd���^hb�O�i%p3M�\�O�ym���'X�d�X� �D9#��$ "1DY�Xx@Tǈs~�P𹌪��k������O���:���� �����l:�Q�X��N��Y�Iټ�G��o~M6��!�A� {0�Q�JQP�����4��Gvغ���,2�M��G��V���%�����='p=P ��4���d�a��
�{6����]Ɏ�DSrϧn����;��Ape�I�Np������ˬd#��x��4Y��B�R(i�a��_8$��?�V T=�3 �b��2{)�χ��ƙsŦ�D�yݪŲq�*�J�t����L�!�{��n~Q|f�Y� �j#P�رCv�V�h��A<uƁ=o<p�\g��� ���FMb$�@��*B�� �N�����F�8�M������6����>�מXiL)��4�"��Sc�a�
����oe%�;�'��CGYK�n,��ٌ<��#2����e�ʆ��K��E�"���R��67[C�(5h�@�y�չ�u�� ��Z��-H����j2-cEx��+䱗ߕ?��$��c������X�y�R�s��;>�hԪ2���iX��diR��a �8��Ha���ظ,a��U�T@�� ��6�����*A�����87�\G��b�k�������o��s��d�K���_�T���Rd����A��/�!�����F���)��0ɢ.����杽
���;D5�,;�:*�%�X�q��Л���/98_P#D9%�E%5,�(ȁ!x���X�J^:9��Q_WƇw����� ���׾$��\�tgϾ*�I�r+E	�.��tҪb���-��0�P2�0���?"������w�J-�%E�i'wjb\�1t��%jA�!9ǵ�*��\*�7^��9�Ma������bn�=vQ���]��;���|m}�k�7�(T�DvQ[�]�C9�̛�≀���{!�'��Ue�hMN@r*"
���*Z�c�����m�u~�� �z��::I� acC��������+Im��,@4d
��D52��# �G�i}]5����%=�}2���r�";�%9��Lwl�6�i%�t����"3��уpV\��w,���-�$k���q�Yk��;�C�>�G:���|ԩ�^J7%��oOi��	I��%UE���m	h F�r��^�v5�q�������8�m^+@�2D�� �b �.��,�{S�� ���b�Z�+069&G!I�{]��rE� �����۱\��n��8?^C�c�����a���^�q�R%}j΃(�F75"0��sn��f� �:Y�������P��[G����KDM����L�>��U�ݔ���W����O��f�:��g~�_?|���W��q"t�B)�	3r������%�l)�Rx2)\��S�X>*�Vo�{L�/���Ti��50rAM��ą��O?y��/?�-�)�rQ�n(P-!�ƦD��V!X:Qx5xL��ܴa�e�\Ǥ�y擎>���a�LdA2���g���G@��ĥ �6Ԟlu4+*1Al��
��ƃ5p�`��P�~���j�PV>���LU�tʤ�#�Mu L�~��F<[���Gy`�e�����9	�J�T��(��( ���r�u�e��Z"O!lV�((����o��o�������K/��+W���zXX�e�l���A���K�#N�I�6�YW�@)�K� �NV���`
' ������BPߙ�|���+l�|2O��iL���'�K��h@6̚W��dg�%���eŪU��c��/��W_�4����^#7 �/�224Stq�{����˽_��z<��Ȉ���y��7�H��m� �Ng 
X':V�j�{%I�0hA�ڶv��/�諲aa
����QX�rʼ�S�R+�6��e�Kۤ��ri�i`���ڟ��?���܃�/�`�c��uW�ds�%��܏��o�7p�NQ^J���o���뵼E�9�,n"��ͣV�y�;n�N�x�m
��ZX�1|��dM�1�\�V�;�B�>��Ƚf����c����xMKl� �N�I����9�9L��� w ���4)��Z��Ԩl^�L�ݴ:�&�1������ 9�#$K`��päa��⋤}(��c��5yHYw.�ƭ���lb�7h-�@� �͇��N�Z�,�'F2�o�(GF��I���hA*S�Y�p��V�@����:�J�w�X�#jV���)QZ�.����j���� �QxP������:6<"?��Z�$�-Y�T	q�~�hǔ&��$�m�Ŝ���H)E�����f�F*�|ko/<c�%C-���@�� 6a]�$R"1�0s���y��n�k�-�d{�k{wWsq�LȵX�'dW�M{����_��_V�z���;��Ǟx@�G�hX���(��]��:�]�.��1�r`������&�7n�������PQ-�ӿ��$Fnx��� ���j��cW�RX}t��W M��wn��;_��h�Fr*#�Uro��m#��Gӣ��X����U�^��&���j���G姏<+�0e��c�0y����s+���J`=���_�| �E`���E�b��~�ix���R����d#���)���U(K��,�u]uי;������zDq����4�2��?����'��ؔ$�k�'k�&��C�i��D��RVn��y��]��[�Ë���[�p�<vX~xX��kx ���63��})�[�)��w��;��T�R�3iB�kV�j�����>���6 k����z�elx�O,��0ZR�7">��ڛ��6$������L�+�=��0��dU�_�-���oȂ�}%I!OZ@]]½I̫'{\��*'��9��ۮ��(���O�c�Kʵ�*��s��I�z�$\��f�^qo_�$����3Nt/�������B�_&�`�w������8���1>|J�+��5�'OH��`�^�aHp�?��3����-��������	I��{����>#���*����8�iy �wn��P=��뇰�����՗_������������jx��G`���5�*�-3��x�j��c%�Μ2�a�f&�k	�������7M4h��O�H�t�`:�J�r�Zn�ј	� iX��������G$ڻ��j��s���.S|[�.L�P���_?-�� ��'�PX���Kى8QH�ό��+���r�ףg�,�4/��Dl3ǜsS����mJ�Z�@8n���q3��s?�����/�$ �KvC��Ҁ��Cta";��x�
�T�aV=Љ �{PFs�;���pm�{�rp�9��AD
�AL�n�ܜ^o4��6�K�d
�_�a��R��8Ȱ�a�J�մ����`�o��_8�W8��P�� ���a924�ő�"r��?t`X��1�kh������c�#V�I�F�+�=X���F䶝[�7���#g�jt�a��ttJڽ���� Z����;a���l`�s�B��ćj�u6�5%jsVF�T����\[T�!�_i��Y'�ψ��=������3J��:��sB�9 �	$�L0+��eIc�ؚ�e[�]K3�6�=�vm[���{$YɒE&�b�Id� rnt@�P����{���������P]���������>��[�b���E�������+C    IDAT|��#�]8ۨ����jm�a�	+CU[��N` �:=6���͚=���7�eU(�e �b�47��g�X�N4z�Bl�O��{�V�7Ib�q�#�v}��޹m;��������6y�T�� ܻw�m����ޟ�
�
��QC[X��Lغ�MWγ��?m��w���W�u�{z�l9vp�O~*�LԳ+-S��
a���� �~�,�ɗ��~��)k2��&�|�<W^F�POvr���6��oj���&��X��K�X�!�0D�R��#z(媤�"���l@�q�*����l��� ��Z�n�D��3��F�ˡ��A���>{e�n,�6�q�E@����[ u���ֈgW^��+:B� [K�`��%��ߝ�h�Z��,��۷�=�`�ۧ�����?:2݁D�[�A�ix��P_�~}N�믧-}9Q�!���8O�DAH!�yR�Y�~u��R��^�=4�7Ӑ�e�I�Ǡ#�Mɢ��p���g�c`�i����j����=���)j�e�j�'���b��	K�a����Sp���ع}�mߺ����^y啶䊥�}C���)Y��9��֤����s!�D(2�wU�ZU���a���a�Hƺ�x;b����ȼ�,��-���W��O^�+P��a 	�}$V�����u0��~��'Cb��/ۜ�sl��lْe�����_U9�����^Tjp���o�?��֢D��@��L��HnT�_����i3< mo��l�Ex�;�V�����>���bc+�����'�������3�.�|.��U�:��'��
P#��Y�c��$��_�8}�NM��aRֿ��_�o��sm�����aZ-�����q�֖�<��Jh!g#٧��@I[�((%g�4�D���X.��e%��ϝI�k��!2"H�w�Nuv���'��wv۞C��(���85iCoX�7t��y�����ũ ]����>�l��j�Y�
�G4xw���l'��wr���>JK}{ ��dR��-�Sq�B�h�`]W���V~�>�)J��}97%w �9:.]�w��4EI�U�(5(�id1w���v�k:� ��֧?��Awg��9�Fk�h��K�?	ㆻ����y��Y�214���^~�5;r䘯+M���u4m�T������I*{M�1�H�>��J5�<w𚏼Qä)�OL�8�Hv�~�>�k��i�j����a)��������a�MHd���+��oF���0c?�O�
�}�Gu�9�5�E���6��/Mr2��u���(�<S;��U��ZO��iq<u��jj�<)���R{��	x��X�k`UVMr�}��^{j*嗯�F��m����RTdmG����N���L8tj����P�N1�($��O�$Nj����m9`��w�&�eq$�=b]�0�/�@�<�>�ظ���4!yA�Y��a�F$�	jZE�!�����-)u�Zj��l:�����O��EH�����s%5-�}�*@oT}}���S[]m���Εaιk�O�o�^�P��{�2���0v���'�q���Q�U)�uA�H/�/W�I���)`Ս�g�e�>���H
�p7��Kypˍ�K(Q%�{�L�N>c�o���d�u�v��$;c�ɤ۷���� !SR3���!k�L>���/�g��3�"���g�8��<�k(�s���3r]b�t���\�u(u���|.T@xV�䚪�n�������WZ*�tz��VE����1HMM��Ԯ��j�H$?�.a�bMQxF�r�;�+�NO����*-��P����;k���������������?�㝀o�DD&���*.�q���K�2��r�7��B1������������7Ƶ7ZӠu�o��X"�1����_���D �X��ϑ�^c�j��3V�۔�j���<�VM���4( t�֬�x:;Y�ѽ��) _T������,��߀�������=���g"-�꺼�
%�d��@�\�;}m���ٟ������ZoA�3Z�T�!#�)�(�KW�H��?P��-T@a8�~����W/S�l T5���dIs���P�.`��J?rv*8Wc��U�ty%�na�=A�s���[����ft��Yf%#���'�8�A�.zV"
�:���m4���$*�g�*"�H5�b���pŬz�e�<RqZ�D��]�"�h?��n�0��BaMɳɤ(ZXcUk�1J�4��8Ӷ8�v��L���t���n�������Mx3��S��|�!��O]�l��.��߳�rZ_�:Y���������7.�I4oі�X�e�
2E��z�('�OC��Q��z*�ޖ���>;M=�a6��0�W%	2�Xy�[\"�[�J�D���ؗ���'cU��Lc����L�ݞy�9knmq�z��]���v ��f�����:�r��x/i8`�
>�f��U�`��u�����͎ĕUJ �T���#4��Ds�8��OE�qk�����������.c;P�#&�L:���F_瞐Ք�j�6$��O�ID~q�P��<]o?ȓ���0���J�u�_v�QAv��,�9��fU7K�A��J��0��Z� 1�_*pR�P�[X��m����;/��T�w�*pT�B0Q��"}
�xJ��P�T�.
�&��'��NLg~Yg��TJ:�`+Ʋ��W*;��ɖ�!�t1��Z������yJy�����{oY�gɘ����i%'�݇�8��8!��NZ2V�_�g�T�qp}qG�����1.y:�eH\P��;s��t~`�T��5V�jކ�ۋ��F�Y�1$/�pa��&�ܴ��� �g�B+�r�
`�N5�$�0u4ƁNY~�u�=v͂ixOt�.=�{����{��Ѕ*ܱ�׽�EuF`=��WB��J��fh�}GeP�ޓ}�h5*���) ��8"H9�$��#�0���v{=2B1dwE�2��5�O�o���㖍��{^WDL$*]�EC�49DF��� }�jm��́�$�R���[�Fy�	I���:�꺋�Ѧ��S��j�z�X����?�`x֮��άzP����ϵ>Ͻ��BAVXզ��Z8T�P�*����V������ �����K��
�8O$_j��K�% sfA��o2	��a���k�}�#+��xF�f�{�(?��$�i/q�{��v�/w>���B?�1���$	R�X=Wp��ᲆ��^ɿ+p�Rm/�`w}_5ٻ�������1��g �u�w���o���4�ÃX.���u&����+����*���o�C mW41�y�PM���� �@j�	 <y�2��F̌���}��g�*r	���� �G}�J2����]�N{a��L��Z��l)ɬZ0Ӿ�ٻm��I����Kf��|��32	�=�~�;�h�8�>�R ]��f[��O}�^~s7�Vk7a["��O��N)��o�c�����z�1SL����B����,���:T�h�`�V��@���'t�*�Ը.����ݴj�Mg��7��=:�8n!Q��4�_J`��Խ��L&%1ɞ�'1�������*�Z�JXľ�Cƚ���P`���橮dAKiJ����ٛ�n_���d�d�=�D���x���suX��n-��2x��VR"!��e�=඙r8楆�*�R �ق�3�Cc|����s��N�+��OdR�5m�,D#*V ��ȯ���uִ��)���1�@��;;;m���~�K@�	��&1�
]z�e��1ӂ�}������3f�ٲ��O�lv����Q_0X�i���i� $ьD6'�
�Vd��H�>Y/��e���ř	�*x���C�@YK�Q�*9+�K��Š�;����HCTx0:b���$)x���
ʴ��7�f�/1PX���Wj�ȸ��#BI��D��s��;=��Td��:����-m	�v1&A��n�}n��v���V�`�K*�霔��S�~��ă.1����r�����^�E&Z����=��&�`56�p{�������/���c4��vj!HJ���n�V�0u���o4�&��--�}�֫��ң3���G��Tf�ڳ��K�zm����TDĴ�`��l%kmr(���xS�V|g_ؗ�W��p���M�I*C*3U�|r�:��s@z�k�
Q}�i���)J��N2���ش~��@����l�N��VWW��hX�<e`MH���+P9q\�h�Y�ڣSI�?o�W��lE���\�(P��y0[��[o��� @��Pv��n�M�v�-7���M2�^�ys��R��u�*�*�`�ŗ_��n��M6��2��M��Ǝ;jw�q���qF�/���}5u�8~OA��-[��n�Ƨ���^sV�7�`��V�'^�f-���%��Z�g@:�C�Ux��0>�'>�����*���o��0f���V�Pҙ�;�{��‬�q���Q�;��G��|��grl����[9�E3Ox #�c�:|�%���&(�%��`�ϗ����>�I�b�<�Q�ޔ�����Z�iTSJ�·�DL	�:l��l����m#Kj&1O��  	���A<�$���2�s�����ݣ	ńs�&����S��C[h�;w$)jd�g�ٍ+R��`�c� S�W՞��W�α�r9��,��|~,"���RkO�qڑvm��5�uI��Bn?n��n�K���>EH:��ܮ^0�C9P���8D-u��}Vό�ysf��r2���׺Q��ܹ�ϟc3*�*�H�Z�����6{�����/�I�?��� kc{��<x��.&YP��w�S��G6c=�
d�V�	Pr��R�Z���/���;��B�W���Jݪ�@�K_���8��sSj�7��d'�ڃ�g}
��\��x�i� _m+V^�ldj��Ǐ��_}���p�M�R�%�S;ӡ#�����0%�j��O=���ƈc�2�EȊ'��>t�{6?���6{=ksk�9��S~��ۆ��; ��3v��M�gʴÜh���?�aȩ��X]t����y�~�ǚ�l����
�"e{V����>�oU^����y~pP�F|�/��1���s�:�Qq��d��r�v�ᲇ� �����f5	�ןa0L5���}�M�����)n/� �T4 �2p��4MG�W��8��xs�^ٴٞC��DkOZƨR(p�?�/�
��}� ֿ��'�Ekn���XG��.W�QI���Ģh>�C����ܥ�ri
7�
�^�f�T����.Vf(���;ȻO�a�d��fs��/@皂�������`s��d+mˡF��\ VO(���$���~�K����X� _4���p�:6J�<�v����������kVc���"C�=��+v���r�ח!��2��ֶm>��Kv�]w�Bھ��UD�z�����؋o��PM�*�� ���3V���sTu��gm�ߵ'|`Pϣ׮����R!��cE���ǋN"�_�>&� P����5_b�"H��l;�d�#�	p��ؓOۼy�lŊ��
��>��
������,[ղ��
0��n�����?�͚;�V���U�5Ԑw�~Ƕo�j7�!O�H���;���7֋�w����j�ocA��ٗm7����pb@���W�s�T�g���U'�'�,g��hn�W]&��*�*8��̕F�6���M�9~�X�u}�;��1��v�Cd�Bm[3�5w;�W�{�N 1X�3�"�?\B9�]�È���P�	�wΞ>ŮY����e?oF�	R�2y&���G�(4w�Lq�^}c���{ ��/)kh� �ڇn�-p�����)�����}��cf��|�6�L��8`=ۍd%X�r��ы�l�&��8	X�2P�5��F�Iѹ~�,[:�	V��^k���5�V��y<.%�� Y�3��{�����Í����7�E�#`��U�X]���Vi��S��s�\E=�  +��Te�>�͜6�n��*KK�&�����&��s/ن�o�UsfQ��^e��y���������6�iH��D�8��'��_o���������㷙�~���k��  {^���S�L�Ẫ.
��*��Z�:Z1j)��3����0����Og�	�6w�g��|g��C9a���ƣ^BslUcu*	NTcU�9s�L�E@�5�TEM����y
��rO�-�|��f�� �+By�O�T��|~ ��Μn�Ff&w3��J2��"�(�A�P�����KO�#.���`1����hW*�T+Ҍ�D\*1�,���������3�{N;����9��Ew��Ӵ���;]�݇,Qx@�&G$2H�^�(Bї��`%<�Hn�5X]^lS'�2�q�-�3��Ϟ�J=�wo�;	Ў�D�s�>�l�Z(A��N�Q�*F�Q�="0��D���<�^�`zpRY�O~��|nL`��/�扦�����e�"鳜��OԜ+��:(�+�[�>'U!ٜ�� nUq�ݼb�-�^�SwD�X���H���z.5�f4�@����{��}�1�-�ho�M��UQ���l�?~�5���*��ĕX�1z�zy
��ƚ=�ԯ� ����}x�e��w�ў|�E���W/���f��bV���>����V[Lf�6�"��J+�X��zP�Z/���U.HN�
�mƫ
��l�:
2��s��s��3V	CB].|�QcU�?�Z9�� ��j�u�A��E|�B �@W�u%�m[홍�z_�+��/2�)P��7��i��(����"�V���^V-\j^�z���&���1g�q�WC&���O���������I�$a�w	%�w�+=��pR���\o3�Xm�����R:@F���K?��Zt2.r���s߳��;b�7�:{��Z�uW�B��n��y�8�� vP���J��tTO��0�7RÅ�/���o]w̿���Ŋ",�Nߧ��ݣ
T��D�2���3�Z�*ߤ�@����V�(����r�#��:&�֒&�7]A�\��)�RvZD�j�+�b�;E�1����CkXx�ZS�5p���7Rc��e�C��Wi5C���щI3���e��6�H kS���g�� ���;�j��j�*b=+/�%l��BүYG%��Ih�CL$h��m�[ۈ�����~��)��H�X�Vrp�0����Ǟ�و_��z%�R6Qdk{�[��q�Z[�|
�&�4P�Pw{����{���>[�x���4�)H��=����mT1�Z���6�y ��JӠ�>�n[k��j[��<�쳌'lv�P��m.u�ZQ]ń�z�ߖ���;��!>V�۪>�yGC�x�D�G���˔���j��w^��nZ:��6�H�ר����O����T��:����&rR%P�z.�?������.�{^�@���-�|�>����Uس�v���XiD������H��ߗ��5�C���)^�i�`r^��,�f� ��+�j���ϖ�-�V�f>W�V�����J��=*�-7��q1[����u�@R�m}���Dc��:a�����h�-�欷����r^�BK������Jg�GES_�-QY?I�������0�]m_��Z���+�����Z�3�v�u��zm��^��+����}��}������p֩����_>3�x��xc���_��+ug&��Я�况��E�$s�RY�%T��Q�j��Tp14������<q�Dn��GB��u��B.`ՠU�ɝ��<�5֎�Zی�f4,�&�X?�Tp/emZu�-����R�V*x���m�h�r�3k�l��W��&+ٵg�]�h�M�e�,&�����g����U1̀NU��˨�5w�m��S6T�o)@uR�>w���ּȣX�8C��j���qɇ|[ղ�ܶ�J����G�k����?p���ت��
�U�V�o����J=���c� 6B�y���s���O~Ѱ�Ww�Ww0�S�=�M��2t��\��#�?v<�a�3��?w���P�(�X��޳��a%uVdB�zV�=� 2 ���Y�f園�?/==    IDATO��=�9�Vى�FtU�������
o���t6K`�W�@9�@�d�J��70l�V�:ܠO~�������n}���F�
��-��P�@ߧ�<�r#P�5n�Ak������0I�_,�ƌjN���\$k7�p&�*$5�34�8��S��O_>��(��; �"	��S�>ԼBs��㵘P�����$^�j�t�mT}PM���;�|�=���ٗ��r�ǥ�����`���~K'�39�R:E$U�nd�a/A���T�[�� B@��Mخ5#�@0�������A�ӿ��\�$�.�ou�(!T�r�QĪ@z����e�R�dKh W�"E_ZG��ʦ̷�y+,=< �H�<��+�cq�9�>�����G�y�R��IB���P��XخZ2��,���-�õ��o�'�%,��a��e|��A@�
V�ֳQ������av�(Belw�u�=���@���o�cϼ�ӊ'L����?�UgP�>2j�܀58D��	G��ʠ�Ү����̪�9F8u��%٥�`K�.u��9r䈷%��-�1
�hN�6�1s���Z�>��O����;���o/���+�k�� �*u�"���#�%�5�$Z��ln ��:֔��b�������-^ޫNV[}�"'Z���A�!p��)�!��D-���s�^N�(-�/���f
�[�]^��ʆ5����^��=k��
X]�0�^����Rd�VE<��6
��v���x%�p�3��@��׊��W̨� b��>�[Kf#E��ݻ�=Ԍ碃/%�ƭ�u nv-j�����pg��m��������rMJ�J�Ƿ������9�u�$��ĤQ�ˮ�#�U(�h�f�h2G)��kZ�K1�жԋH�i�/U'4��ng*�Z���6\5Jtҹ">J���^�^���k}Fc��Ls�.�35��Dm*�ä�:;vx���4� �!3*� �{Zީ&y޴�F�?���0~����؅�t���=��5(a�+l���k�܎j�V_�u��<cM2�|�^��@���o�gJɪ*�Xkt�:�8+���a`�u������o�/�+���Y%��2��hlz�7�m�vD<�h���B*AT���<V���>@rT�һ����������[8s^[DH�o)�������ji�c>��ĉ��֫q�e���*M���A*��z=��@�R��6��{Ȼ7����R,W]c����U�	����K��O�l��<z�;J�h[�&ʹ7<�3���_+@%��k��bj��uJq�'��[��/`Ջt��.J���:��U���Xua�Xǩ��53��jsRvǚ֐�����iI�����5.=���s����! T8?r��jl��ꉶ�p���u���Ck!qE�`��#�hۿ�kuU����&�Q�- %KJq�����TT͎�$@�ϫ"I�2(N�|��4�y��͐e�LE�:(+&����,[=ɺ����Ha,��GX}���P�>�I� �G�s���v��eV���!�O=���؛�W���*��f1���!9��B�DB��8�1���r����)���^�j��n��!��lf(F+��D�`)��3_�Ay�����$�*^�k6Fk�ڵ kQ�I�=
5V Q�,_y�Y���{�Ͼ�gv��Q �{���2��k�yCf�� H��(!��rD!`��E�S�I�U����L;ܟ}�O�C��Z��UͶ�����n����O�� 
n2��v뇅�*��UuV:!�X3g� I��'h����m�|߬�E�Ll|0���A��j���� L���s��xכ�A���r+��i��zr��L�eW�\*�R9�7<U05��#c��m�yI ��N�Jm3�\�
7����M�@AW�(I��`1�M��f�HMH�/���|�X���!Eޞ�G��e#��-v*M���֐�������n��Co������	|�}��I�$�륀Kݨ,�L�uA��&u�����L�ueqk!�@��5ֆ�T�ڱ�z�K��ika`�C (`U=NԺZ:*e;���:����ڵs갘���{T_K�(5�����i��	&�0�h��:�P��L"8>9v]�G�������!���q�ZJN�cF����Y0���}��w]�*Ò(�
jаf�E���/Ͼ�X��i�q�*��Xq]�
���55f�N}��wv�j��_���z�N�Jp�z�L7�ߺ�͉%~NoATp�(#e�daǎ����/2�u��zNun(�����j��,��
���M�,^>�w闄!az�oOe�L�Q���q:�A�8�'�y��&�%W_���J������SM�g-�uw�$7�4l��5^�"���E�+c��
~��/9�:	*�	t��υ7�G�����Viz�h!��J�_�m�3����Y<r�	���V5�w�i`P��q)�UoM�8m�&L1�41������{����&��V~���Ŧ��1�vZ)�NE1�L�]��5Fs�Ϩ�K.AM��6ED���j������z}ՇW�0�uȰ2�j3�,���IV�`��<M�?�knxObxR���Uh����޷:Dvp˵+�]j�dA5�o"��ٿ��}�$�h�Ql@�-1	�7\���\gn�8��W�!U�jl�(ToŸ��!^b-=�y����;���n�	\Qآ��F�a�˱��g=���y`��K��j��?�X+�־q�^NY_���m;��j�*w�������9�9�� ~=���)p޷o��
��X�W2x�ч�.Е� %�҉.^�L���}4Q%����㾕q>�O����
�lHk�\�z���އY�R����&ʞчk�,�Z8=@�\�XJ'�26<�������q�U ���q�x���.����*�lT�i��[��*��j�Ʊq�A<��(�T]��X9|� �H-p���Rs/�/6�W�u��̚"�k�R�e(�Ztcu��0������
V�M�5���k����#����n���n���7-,���>!&A	=��js
V6���Otq�qCը>̵��cl�C�.O��o��IlQH������K
�����1���C��k!F�_����Ƨ��?e'�}�A̸+�w�lH�<�S�+���A��R��EMl���҃�,�t@�Lc��D��3Hm)p�#\�����z�3�fl`�5N����6!{�]��������8�^�U�ۤ�v(;l�$�(<0�{9���0���o�A(f�V�C��s�`j�M����5W�~Cm�;t�����S0Y �t>�r� w���q]����2�^�5뮷�6�c]�u[��ݶ��>G'`�C��)`����%��}�q��{�Jv�v��.�m�X5�f��Hh}����z��J�) ����[F�-&#h%3*���?u���C���*��ᶵQQM�\)x�H=�}�w�4�6�r1���~��b�P���Pg@��m���ؔ)�_�=뤞��έ`�Hn9k��v��Bpk[@��-��{�t����@�Z���:2�A^� v�i�NV{��oC-p�N.���o�W���Vcu`=�-�i����Q;"��ڱV=b�V�5�X�|r��@� 4�Օeܔ6v���72Y1�H):̂IAAݴt���a��A���0s2����r"'�w�=�3��Ae�N�k~����v����n5�N?tT�E(����j.vi~h+p%�z�t����� ���ӽ�H$Q$;��oM��VM`�׀�>Ҋ�q_����o��^�5�*,<}=F�A�(6�/��V�?����(�s�'��-�	u��f��^��iM���GxH��6}�x"�b^{밴��:����>�b,�+Ơ�5I�Z��/� �,+fXa=�^�����$zNYr�U�VN�	Kn��p���cl���z2�c��5L<�$1�
��E`�h�O���9}�V2�(E����<���_@�f��kq�+9����Z>w�-�Vm���U��a-�yg����3hh�O�:�Iۆ,/���/~�?jԠgR���/-^��Z�%v�k�Z�X�(T%���?]/���:�(��zN�; i���pU�(S���:���L���PԾ��({c���s�S��}��
 :>�Zd����\�43QӰI}�&J��s��H�i"*�2�l�{�����ZeU�}�O�nӦN���󿂀N	���|Z������'{p����wvӌB�7c����!�t�f��3���8�7�ڃROwO��<��o��Ɓ,���FX������RSݰ0���T����k`�ÆS��F��SJ��9�m��I/\�($vp�->��h&�����ڼ�S���Y�D��m���h.��V^4{���M�ptNЈo�D2k��֮��zwpI�)��������ڈ���&�K3f��T��qx��*!R<a��N9�����m���!� �>��"�(��$���u��7��Fk�&T�wꠥ(λg%"QC�j42�����2�(ţ��R|=#`M��������Y����ֵ�u2V�$��EGb�`D���="��:�� ��-�\�R�F 5�ĭH34y��h���T�
�.�����^f���+�XuPr�r��YjEUm��Q��p�X�&IkB�0�CWB2k���Pm�.r˵�즕��A"�j��lz�����W����gd�i⁓x�=����Շ��-����釬s��^�v�^۾)+��U�/	B �b/���~{p�M��"P��T�(TX��BI��${,������ːR���a��_�ǀ����|
�rA5�<��ℤ�lCB��uFj�]���ɊkY�����3�j������g���[o�a?��O|Ġ�0I���}8O}Bo|��6a-?x�X�}87����`%(�0[焄NY9JͮsE�:�94�"�����?��G�}��V5�|��p�tu�yC�f��t�ɰc)����/�7�֭�@�a�(��8�롢�>p�g{�J�E��6o2֌?��&�K*8V9���>;*�,�l�����D|�&t�yT���E@"����;�SW8r���=�ت��1����@�Lٗi�����Bw���1cљ�7��' Q��\��D�C,�7���˓�:!?�͜q*I������:2r�u��p ���U=��A��OE�i��˝�Vں%�\�WQ��ӫ/�l?����������dM�f���1�ˋ��^�e:�(���z�g~�"^�q�^߱cx�4�)���R���� ��+�^ik}���{�1�' �d[ߧ�I�({��X����F����q���?�R��(�9����Er�����xG�!��Ag�qv`=do!^F��P�`���9�n߾վ���Ҷ����TW��5��3��h-Y��&OE�L�c���VXg/9?`%c�Y�}��o���mN�X/�F�V���{�f���q��u �=L�e��O2q}��d�E+�<K�Z8�j�z���	��N�����m���dbN�k��XR ��8�M����X���� ��b���H�6�q��íLP��e�=Ų�ἥ��ch� ���Ύ���^���'�ʕXK`������F
�CN>�-I}_��B�]i淣S�N�����Ê��ކ"F!�P��g*X�`+T��*X��bT����i��֛[��'t�v�ٚ%���sp��[�֎-���'�p1��H�%#O2'+3)�8���y����8{ݱ�>{�/[{�כޱ�6�򆩗5���"	�2g:���LTN���I���g�ȼ�Ώ(9�<ƹw&Qم^��z�'�1crY*��ΰP�gTg����`����9�A$���RM)��惶�Wd��L�6�������t��c���������W�,ǌ�ȕ�V����vwwڶ]o3�a�*�XW��;��X�E_
`�5�b�G��?h��������� &�kȠ�%�*�uʦжz#}u��V��zl���E=F�s[W�g����ADN*|�����9��|�z`�a*�p�jY�2ID|1���,�q������kli��6l{\�4X���[��1F���f �^6�"�K=rb�d%��|��&_+�=�����V^q3D��i�HCj�@C{_/�F��d�4B]�B�W���6c�'P����R���R�g��\����,�LG�-�?���6�u��t����ۦ�^v+J�3]�� k��������V��ʅ�Ԑ5H{��U������C�v�s�z.]�kz/�����ڿ���v�R#`ƢP�Ś_,-HAT�{�5M�ljג
`�ߙ�{��z
�Uu|���������"6L�N�r�� Q ���F,1��0�0�rж��v|��N���:�<<�ߵ���D<�T;G�����u��+l��	��Ψ����}�cf�w��_=r"[|��IGPS�UT�.DP[��s�Yd�N�pH��\��}���D�v7ی��r�[�p��}�L=�+�&e�2H�Ֆ�%��$Z�e[a�5R�}D�?��I��G�m$�m?4��!��z/�(���$-5�E�!�ľc���͐o��eTr	���>�4����z�#_O��&��������ك6�j���TS��B�3
��ѓh��������]��j�����c�ń}" U�����K�T��P�RWS��̬ӟ?�J6*= A�(��Q�	����=�����֫�����r��#T�v����4��XuI�A�u��~��(%�������PJ�"85�V�B�+#�����J`�7�\���P�r+�X���������AS��#���z��<��f���<y���?�w��X����"�r�f\g��[)���Tp�҅d�P�OB?8�V�������Uh�M�є_Tp���jW�Usu*X�~�	���<{R��^<�fM��*��A��y�6%)��)8�f_����_O�c"^�#�Y��nR>cto���=�KU�_�w2P�>g���j�H�.��m�0�*�^�),���LÂ��%�jUy1�� |�X��Ǭ4f���cL��e�(�!�� ��(=Խ����*kJ� �֠J��L��X/2�-��������aZ�,�p��6�ۯ[a�.���(AV[�������~�)��d#��ퟰ�t�{�������E[�'�{MH����퓿�W05�g�|�^xs-o�\�5V��JO��*kx��5V�2e�r]*�`����_o&��6O��kx!�z��~Ve��M�R0@�:�1Ns�3�\��I.���=�8/�,��X���� V2�I&�}�lޜ��k�����QT�j�[wb�A��b�"��/�\9��ƿ����
Lc_S9�3'�`���`�Wm8���`���C_͈��uUO�S��v���,&��i^$���}���O�y��C�o� }��X��Ǫ�^cL�_@9��/�@���������Y5b<0����SP�r�Ia�%��V
�[:�x��҄�f�n�(�_�B�C-�$�KHb��b��ď	�A��ڮ��IV�kt�M��@��`�(��_<�h�z����kא��8 o��^��������S^,�pA�6�X�K�M�b�d�X�q��V/�;�Y��r-D-�k��b?��XK��(Ƀj�7z�֐K�:W�J�t۝�������X�}k����ۗu����x=���+W��z�Z͠�L�u�*o\,A���ߗD����laϫ�_-7:����<�*2e(���J�(� �J�W����<��"����?Bz��/}�O�����m��5V�����Μ�j���˝
V�U�%�X��,��w�<��ӦW>	�*c=�+�Re�c�9j�%�a��T^Ze�]P�E ��$L��f1yF�;��a�&�ڵ+�?f1�HVydb���^P�AWW�5���1+����'2�q� 8Y���e�{_��� Q�� ��+eb�4�g�(f����U'�n�7���3\Ym�/O�||1U;m5��c�g�NPc<�_��K5���a���!)Q����e����eܫ�KIϰ����s���"��4� $E�c�&i�i�������BD���r�x&�_�t    IDAT��V2��Z���׼�Fq>C�})�P�T�n#6��v��kX�>��%Q��5K Ӱd=��ib�*�c�R��9\����,�GTp����+��}QW��Ⱦ)�8���CĀM��� �BT��s��*�����c�I����}�S�����&��5׭��o���mD�:�dY5�oƚ?/��X�������/��t�U�����R(f_+����$��٪��I�DA�S(Fv%r�>��ߕ〠�"�v���|�n��[2b.<Ϣ�3/-�@�By��Ӫ�#A+����t�y��U0��
�k�	�?��ڢm���^c��pgt�5��F>�˖^iu�~���e+8BI�n#O��v���TRq�&`FU��'��[�X� �?��GN��~�Xϴu"��n���hn֯(S72���a����a�d�VBT={�[0k�-�5�ԌC�k���f���P(3N�8��e�3%:H�@�$��d�)�ta?�^��eѢ�����dZ�?��f��{A�������\��A~���AR��G�YDz�\��S2���9�LFR�9�R;-"8�y��56CʳU}�ޟL�YT��T�Ԁ��"B������ڔ��F��W���@��
��>�2����>�pp'y��>V]�0�؅M�\�ǊG���cU���ݢ/�ʅ�:Z��9���Kf۬	�-j�5�#^������sO[%��D�+�\���sCmx]=�6o�R[x�5^c=JŦ����\^��i��A��l	C����;RSW�'�(Ï;E��汖$����� ��� ��|�3wt?�����A"	��˾0����G<t�
��ӟc�GB/-6�n���֛t����6���yWL�ZO�̀�X���	X���:u��o��>V%5窱J£�l��EV�P �'�n���
V����B��Ԫgd<D��I�љ!m�s�>��b>�,S��j=x`6Ԕ��6g�D�9�ƪ�Ɗp�Qۍn��_3_eF��(�Ԁ\-�J��X}D(eE����U�=-�^�i<�(I3eիZB�L_@d[��v�/�XiسV��Re��%�����`%5����٫����B����Nyơ @Cz��ߜ��#�E��b��,���������%�(NB�Ri�W9�h���r^tZ1^*8�!�8� "R��6(v��돁��"��o��Ku`
@%^fƆ����k�X���٢*����>m?��O�:�r�d}���HV�R�X���E�|�]��S_��K�ګ��\��7= �Cj`�tNr6Uq���܄?�XF�B�#�'�l& �LV�ӦM��s�L�D!Z��$k�Yld��$����
V�^�<o�<^�b� u�T#��y*K�^�m�1��b�Toi-tp`��c�9-8 ��SYρ��u�#���uҤ���:u���lӦM�	g����Ю���'Ns�%�v����n�S�y��C	����Ĥ���ޝ�T�:��Zo-9��e��\+��P�h��	55��&�ڤ�
��kÚ�*��)�ue�%3

�y�G��kNP�_�=>E �0��T�����B5�aP��?��geh�0-B�;ġ	`���%���jr`&K0ee���0�2�J	��&�\�^"�Lq���:�2}�Z��Sd�Y�S3���p%_n��x��Q��4�,oz�ղ"\u����YG�d[�6E���%j@4f��^��JI�U>�n̙ �2�l��
f���T�g<g�X��i��YQɅk)*�����5�l��V�׆"�� 4e/<��=���ypZ5�Y������m��R�X��CT��5D��u���e��|�f��$�{^swBmR%�0��� ֞&L"س2�`o��o}�*-_�܁F�y����
F=SY<��N<���-��z(G���d�����^���`��o6x/�f_9}�S0�`Z�z� �`q��f��u��?���' ^R�U�%�'i�
�#�{&�HM�4�ݿǶly�^|�5����{����s��3+����y�eOFHcq�y%��.�����^��i?�IqQ(�,��k*��&��j�30��gN�𤌃@Y��q�N�&�E��� ��2�W�Qޖi��r�LqM:E���Ȫ��Y�y|BKb��f��0��y��k�8���/�/2�1bBLc�1�w���Г��#j�6^W	^)�Ф2� �,%��_�3\���}0�`�AM��?��:uT���:���~2&�m�5a������;/�X��sk�Љ�2��먪g+@��%7 	�oG��ur/��M�*�"�Ep�\������~鬉�~�<7 ���]۷��� Q����J����!�������:��
�x�/����&��A��B����ֳ
�}l�T=��U&�e�+�cu/ ΋�[7�-�|¾򕯸�ӃRg� 5�3ҹ�5)���-��H����D�)�ܹӾ��oڒ%K�Cߧ?J`6n��#����p��+c�)��YE�ʙ�=+V����`�j��c��M��a���n��>��`S��46f�!!y���5�᝝%�W��Ƨ��̿���{��o~u,k�^5ָ`
��|�_,.�n�n����p�[�FZy���NP��4T���"t5Y���u��V_W�$��<I�~qbN!Ыf2b	��d�IoC���U��H ����|j�]�T��Y����=-c����ZG�ְ}4�W*ͳzK���hj���j.EVᰃ7nS��śwZt���l��V�"?�R&x����u����A�7ծY>�3�U�X"�S�%��[;�J;����K��7c�>DXQ7k�
�������k��0�Xu-X%В�X��3֏�����P���X�H��v댆rgm��榦�擶��7�?�2H��SW��G�
.��|`t�o��
�Pq���|�z7�8pj���S
����3��9� F�
��*`����(d� �A������������|ƾ���A�H���Y����ۛo��$�����K�p�Znݼ���o���p�z;���_���R�<��ϙ�M��A:��x) k_Y ֬�yy�&T��UL�pU0�tp^z�1T� �v����(.TEe��
�z�!J��5ؼLz�Ak�f����Ϸ�:�*��������X/G`�'La��m�:��^�O��M��Ӻ�p�������8�����ՠ<��ڊ��y�a��TQ��F���.
Rm5yPe�����e�A�oS�����5kU�H��U�{�/g���pN	�J� J�;/�:��,������[>�>�~9vf���q3��H�=�ĳ���l׭\b�x�o�^)F�'�����h��-�z�R���uV��,�M�,`���/�q(�~C������B�ҙT�g����U����|�5�Y���2���+����D�\0�n^������Yg*��c�=��qo����#׾���} �o�d�ץ@U�v�4r��R-Y��V��Ɂu_Kڽ�/w��蹬�w/�R��y�)�K�|>��C"���e�.��
��?����}
�4�U����1���ӕ�^��6H�� k������-o�e�u�����6a�$��Rv�Y��"��6�SC1DE󟪾i�,�6� kFBJ�w�֐�@kgPc�.��m�}͇l�?��Y�����?֝��9��v_����3r�?��i���_=?*�����6�vcΕ�3@������ Z�qŤ��$	@}��!J!���lR�)ܐR�AOC���� �4ũ;~�`��A!��e�a���jx���1Xlz�pP�+Z����
��"��T�mz�����q�t�h�u��ۧnX� �V~�GE���K�#�~	�甭�r��}�2+�a���P�U��Z#�W-[hܼۺ&�����zK��~��ykC��'�
�F�:���X`��P��3�ݿ�2z�R���v���)D�j�=��.Џc�g�������V�Л �+��k�{�|"����3W5�&/Y����d�G�
=�=�ᇖ��7N���ƹ$�W�3)�	V5/����믶��f[����JH�����3�\�o�b�h��8��{ğ�/�G�����K�}ý��/|	�R�=�y�=����X'���t�dl����V��{���܈���_��R_�&8&��@7�`{�������"{k�v��Z[u�j�=s���cG�z�3P����}�=�ߛtgT����_�U�^���}{}��[� �x�m��&`M�Q�^	�i�CZ��h�I�݆^͡����0���5a���������0/؃QƂZ֚s�M�!���,�퉣���)�\(��A?;ບ���?8�zz��IK���:��;Ξ�M��0��[��{���CE>d�Ye�R�q�r�.�,E-�8�W��'a8�/���_��@���������k�d܍'Ȯ#0�����	�e�Id""�
���}KX�: ���O�/�r�cNͲE�Tj� ��^���ۺ5����맠���H�������U8W=t�j+f�J�i��h�ԋք�f{v�R5�{9ߒ~aDt�*C�x��	�d2�ѧF�u����<dW]���8T0�ŝZ؈o����ﵛ�[�޵�\��)t�������]m�e�
���4��w���	3��H���z�(k�jǢd�V�8�{+���߯��1��6܇�^n�X9����V�<��_~�~���!z+f��*:���� ��l�[`�a-�U?~�7�v�}���x���[��]�`g��5��"f���T�K�R
�΅��~w���\(�yيBŒ	H(���b�PA-Q}�\�$�S�n�Q�ý���_������%�k��?��(N��!�h⯏��U��օ�%��a�Z A�X�汦�AD?�h��ꗷ恙�^�2n�}'ڶG��"��9���묥����6��i�m5�]Gk.���E*X�`Ir*f,t��QO�zf���� |&`��Q�%���_�3�.Hfw*MsAS�M飃ߗQ�UQ��g�C�zcE����C EQ��"t,�b�A�^C�&�q��}WϮ|�L XW��yX�
���.K��4`�E<}V�3mDrzR"����V2vݒ9���U��5Hoh��x[�~�����îXo^���jI�k'؉t����g�$nPW_1�>�~��80]F��Y��0�\j��s�h6�z^����[G���뮰kOw�7�}����lÆ;m"��{�	�?��.���C�b/`Ot^��Us�į��~��;�~4_˰qۊ^�a[������G��A���sa��=,�8�A�<�i��HK��5��s	���gVx0��N��q�1@����H8ɌbuX�Sn����{��3gj���8���$4�{��n��i��,����>aϣ.���;.��@�.4�
�Č\��?��x�����u�������P	�Ua&j-�Z��f��NVB���y+����1�٢�'���5��q�峱���	���l�L!��1l�ظX�dVM�[+�L�=)��ƶ�z�폒�v��yx��?��>R�J05i�$����;_N�+\�N��9���\x+B����X���_���`�m��x)S��@�CR�v��ʵ����lU-�)&2s��%�)�������s4p�ªi(��շ���p#6%}�#�פ$���tp\�w��꣙~�`re�(y�)���J����6���b��iN�]���G}}�6g�t������-E�Ѕ��@c�����K=6��m�,�5	�T�Z��6v���v��y��v�=d��j��Ȉ��%@��y���_akπ�n�kULc��� ���޻�Z�C�D_aX��K���l��>�:�����7Zo?��׿?���V��f5x�g?�O_�i�۬V������GX���!��*SQj�P[�+CKâ�6��� C%�C�p�v�� z��V�.��ǣ,b��W��A[v)��*x�C;,\h����D�Ύu��
���Ok��/v���=�P �t�Qe�2����W�Z>��"���S¤�P0 �-��O~�!�p J 6��\��XG��������o�r�(�e4��������{��āUɈz�C�!`���uG�S�Lu��%�#��d�=�X(]�C?�=K�X�&Y3��e `�Ǆ�B�uFe��'��[�| 2�ѷ�l�i�!J�G�!���P�f's���˩�	h����y���^ղ��]*[/�甍�9"/�5?Y	:��:��h�ZY+���*�CI4Fr�(��HI��2&}_�v�5Rd9��e�Z�ЧL5DF��є�"��R���ΘD;Q�j�O�9v
�F����X�o<�����=r�jne0Af8��S,.�fO(�P���Nچ�6uC�Py��Y'��ЩwP�؇�MYLt�}�/����@'ua�[��"{ ַ��w�i5�z�pw8���/�fXF~��w#T�fC�xe���Xed��ﲺ�.X�ed��A5�􅭶�Y� Z�|����	�Nyp�NV�p.����ɉL���n�<����V�U������^}�~�����fN�ߐd�!! Ӡ��R<�yj���gx7}��y��օ���}���΃���>dg��A�{��%p	��j�����N��!e�:s�r��M!V��O�6�R\�R�WU+}D��%No��[��5Z�XX;�z?���W�#�O�G���)�� ���̞� �h�� L�Z3d�����Ug��y�B#��Zjo�~���`��j� ����l�+��0N�)/���կ$�]8�{Xe��߃qT�yD|p�u�e8̪��Wi��@7S�/,wg���D(E2M�.@���j9UU�uW����'
�HmAKH/�L��Q��U� ��:��(i��TaG�8p�@`,�R�[�M��ЗW��n/�vS�?ud�Uѣ�R��*�G�_�r!P�ҍ�A#�7y��rjL��պjX�_+����"s��>���zO��-^�3��J��Y�>���֧|?�a�]�t�bw0��:j�����u�M��9+�J�E"�z`mll�/=��Q��uc�·}��/|�^�ȴ�1g�����=���{����b�YqD�GXuOB��e�A����C1����?܇J���� b�$X�x��K���������%o�IT�q��~b-�\I�g�z��hn��N�}����7�񮽼ue�	��/��V�T�o��5�L A��L"N�[��~F�~	:U3�����2IwE�@V��y��]�?�qH� οA7ta������a2���"�i}�������:�����%�k_z{�D ?6���>F���M�>��������o߾վ��8cRh�utf-`�<�	�r�X56N&�Wn��y�X��U5V5��%�՗s��ذ E4��#�{��� �'{YPP�R���w��^�4<E��2ڴ�?�'L����[��$�k,���{F��� V��>j�1~֍�a��x�v�J|]���l���{�s"r
��4M���]sસ!�(�rq�T���쵶C�l�j9D	�\U�RŒ��0ʷ>h�*��)�P�l� /ϒ�f$|�N5��D �		 4,>��ᰢHz�����/�ކj�9sZ�L��3ݵ�y�Y	﵂�x���6oZ��r��b���'[:���c����V[�pF��3%�c�>o�aݵ^o��%��2۲��뮺�����C'n*��}؎�"�I��2|t�����V�+�5�����䯪u�f�	dV/�c��C3��Z�4��o�a�����=��Xr'K!_R]�:�Z�m|�ߣ�4��nZAn���̗~�v�
{�w��]��;�<��n
t���#c��*�4	�X~
%�X���)g����YϜKb�\�����8�ｈ�|A��3ט���߯�7�y��s�I�pϒyIb����M@�=��g���x��U^�����t�vm����:���	�;������J�P�p
�ңגX��W������[tKC��v�2�R�    IDAT[~�g�XgV=�<VQ�,`����T���v�A E�i�e���	\Bw#�O񧎚�<|1gOc�Ie��LnaݤE�q�k��V���k0��:�j�'�hQ|�e�Ϻ����@e���]�s�����k�P�>
I��/Q�R��&ҧ~�\��7�G|Ϲ	8	�z��@�
�BQ�~�:���"��u�*�z��%;S]��a�W�GJ�^��*tz���#��%� T�+!��x�Ȃ���.��	�׺�6����܋�%��<Ђ�G^P�`���R{'G�2��ՂD8�ٺ1eV�O�| :@ſJ2y)�ɬe���J���b�5miڊ$lʰi��h4g����D��]����`�\>c-Vg���%@��W��kټ�V�n�R��2�2i��d@��z�W}k��Y�)T^�d<��zka�X+4
{�XW�Yk�n�����H��>�Qe���E`�צ0 �tT�^M ��jo;�(�gm�/\!*Ug�%0сh��cO�������5C~;�������y��������* f��5�㭃_)���|=>������L�٦&5�9�f���o�ظ6Fu�X�ł]�|�g��p�s��ևӏ汞�*�C��!jt���aŨF3��na(:S^���-pg4�ۂ�Sm�Dl�wG�nт�-���ĥi���z�J�2�~*Y&�c��s�S`��&�.�G��i ����^������ޓ���)���qR�w���M�Iԩ~�(I�9Ծ
3���r^�G@TO�Lɩ=����X7)>P[���?xCK)�����JePߖ�0U�7h� �YoĖ�c���!��M�*�42	��9Pfӗ�l%�Y;���M�
�ވ$���޴!1V�)�Y�i%}Qr�Q���v	��mK��	�[�ݣ�}ZJv�!$W�+pF@�Z9�����$Í����I��Q��Ӫ���,��_�a�gA�>Z��̥�f���Sce�ՠކSϯ~�3�ˢ�'P���E4�g$���7v=�`Y�>�Ͻ���
&�Q�ק�c٪5�䪵։o�����il�!ؙh ���=�g=;�������FN��C����e�$�;��
ȊYf^��5�P���Kd�,[���s�_ERPI^^�Y%`A�)�CO|$]�
5]����f�#�!�i���:��?�#[0o�S�Vyˏݟ/�6��_a<�"�j��{�:�^<�2��ƿ���cf�w_Fc�r���,ތ(�3�t�����rk{+���B�5 5���N̞km���6s�Dju�n>��7��������-�����>7�ws��+�g8��6�!�]2� \�O��G���M=��=9l��Q��am]��hdZH1�"ͬ��}}yyr�8�ŧ�-w0�x3*廀tq��P�>˜x��{[�X�S�>��|��ϫU���&�$f#^�-�ω��W ښ���
���JA�k������T�lO2ɿ8*X�)P�}�aS�t����7d���0*H��s4����KUg��g�ڈ�~|9I���F� &D�*fS��pD`+ �Ȍ5�7t�q!D���g�z���ޛ����T[�lE0 x�穱~�����*�gbM���Y]PqGz)I�JP��/��S|���5���P���� ��Ǩ�V%�2r� P��+p��|dH�N{�{d���+�G?�_3�o��S���_��|�o�mh�.+q��X����b�n/%�jmƀЅ�-%J�'����ʟN�:ŪϿ�,���l�,d3����d	��,VCk��L����wN�&2�������ޱc���	K'O6�Wƪ��z�U>6N���vU����Xk �_].�Xs�!֨���e�Ѧ�pr8?�ߪd4���6X���@�$��b��f3��
�h�p��jj>n�8��O�Z�~�`��2��#�+�e�ɭ�����pH�n�k����z���}�5�ԙ������$Gp#!yߊ���y{Pr�'F^!kMD1k�d0>��H��nk���MFD&*��"�(GB.s�"28t2�֡2�y�@]�{u��5ɂL0��DP	�N	}�
[�� ��>��km�r���+^*��~��y]�H���|��}�AQܨ�2;��h��J�9t~p@�n�㣛�F`Wut ��g�R�G̝�gݴ�J���T�Rl�����^���_|�� Pe_oʂ�}�z>���=M��KF�����]4{���@���8�=��;��Tb7 �n঴����-�s��r։�Rϯ���Y��７>�߳~��^��\�7w`�	��c�MUsȴh]�v�����2�hX��c ���Q�fxݱ��&E{`~�B>��@��#e^�h�b4���E�M�K+�����Mfl\V��*cU�6�b�_�3��Uc]���>Z�H�XQ��ͷk��y�Xϖ�^V��ش���va)*X�|��`��P�A�`�"c��(4��ܖϝiW��l��Wk�Qjm>�L@�����*����ͯفw�uW8rR��N�'i ����2v�V��^+��{��lI9�N����.�Z[�i'Ouٱ�.�c���U��u���H�j��
��k������qp�բ�,�,�Ë(�y�ꮬA`o����k�苧�_�Z\.|���Ք(�׵��{8]VoW~�f@}�L�b���d� #�yޚ����=��?o��k����ogrO#����ul`���MB���.�J��Es���iu����uHܻ�^x�)W��oQ��q|������<U}OPe �Po(���hz Y7U���qk����X����ki�`�˗[�4���Zz?VyB�b*����Y�%�眨]5�L�j���u�2�����C�_ٌxi�N7O	{"�(s4�e�ܓAuG8cVg[�d�f#���j��>ƀJs���x�{>���{
��:d٣ۗ 68���IM�I?��'~h��al�}��%K�����|�ea��.��.����6*^�^5��ƿ��cQ��%��EᝇQF���/;P���ѐr��+ TQ^�`sh�H7\�ʦ ��lk/���`*� ��[��G��U��C7bΜ9v��u$�h�ᅅ@ޕtʦT���Z�>d\K\.O2��NYļ�4M���N��on����������u�!$�-6��Uĳ�������zu�)!�l�c��w���ȃ�X&:W�R��k��#�TM�D}�P�j��4���\\"���!}gqF�z�*��sÅ!z�����V�
ۊ�j��f����2Y���?�5�3m��yCm飬
I�j��X�*�P���oԓ���N"�jy�3]D}��A�u�YG����8emb-Jt�Q�ܬ�A��Ŋ� ��<�X�����9�V�+PM
`�L�g|��L'����|J��`��>�.Q
h�~s�Lj���Vp������R����T/��I3l�ҕ�RL{B�H���h���6þ��X@p�U��^�Oi".B�����s� �;X�s%�]Q�q� ��d�b�|�y�JT�!ۦ>��,'�*8���n��ޙX'*���&��Y��c���,񒀵��6��y��2��X�:ZY�?pC�U�$`tvtS�����nj�IC�*Z��u�TZg�[u�M��p{?�غ�Z��,��:�e��z��k8��=7+c��{�*�S��F~��B�<AѫqL]�EQQ�D1|��ݎ��fk[;�#��S�x�5f����k � ��&R��!��kz�N��f b�([�4m&E�%�5H���A��z��-�}%�0PÊߥ��HI��L\�AK#&��YY� 87%�I�]��:+����5�uj�k��|F0�b�>[@T�b�A=d��V��3J�������aPS���,�3}4k�#�5RgW&u-�bTO��L[�fj����R���~3gr�]�b	㽨����ۙ�9k�L�5{���4yW9r�֬Y�����ܺu���ׯu�t]ϵi�&��]�b��V�̢����9`�N�5Tډn�!W��~~��W}�ܹs�&[ZUk��؛��Y��.���X\��P]	�	����� �Z/j����ʥ�]Yk�sK�K � (
JFd�|ݳ��������{8���U��]*3�@�jU�K��au$5�_���b� V:��Ǧ�Fۻw�[�F�	X���*8w�[���aZxh�!�������= ֿ��GNd�o~?-�^�9c¤n�����P� ��ɟj����v�D��-k������fk <�Z����}����S�:{p�!K���{ ��*��L�)3�'�PB�"EPD\D��]wW�]�]{�u����H靄 ��63�^�)��s��μ3�3��]^��y��~�=�)�y�T����T��I��N9�4�)qf_@�|X���FMh�j���-1����ʑK�9cI8"�lj��m���Օ�����6"%ؤ>.X�R��u�9tm�e�:���L8?���v�ծ_��>�6X���OT�E	� w��%�o+��M��o�|WW��J�s�ǉ�5ua9-�S^4y	F��,�t��%����X�k���d/$����;ݢ�^k
�81!�z̬c��x�6Y˘v�u���u���v��H��Z"�o5�XS�dl5�<vo�MN�d�v��7��j���ys���i�������SC��ZgO=�s�9a�j��������>;��$��N����@����|�A;�3<:��(!M|��w�IUi'���^��{��H�>}z��.(B�s���ѧ��L�
if)Z�,�O��X�aJ߈{���������p�#!)'�����t"��|�ގ�î�!��� 
��g��TCɦ��C���`�a\Th����Jo�����\a#���S��ݙn�q�tol؄6�����'�tV��	�،�>�[�:*��{��S��
~'�5��HJ�F1V4t�t��9<M�E��G��RO�#�َ\Wy��3m$�_��"�[S�ٖ/C,��/��~#�GK����UϖFm'�61g���duo&���G�=a���2D��:�I��>�R��A D�*dq����l�\S^k[� �l%%��&����V?�|RWɤ���)�d �S�/�3}�eYe�V{�����
8�S�j��v�R{9(�䳮MH"*�<m�`��륩[Q���+m��J�d�EҰx4F(�=�$�ш)�����겼��Jk A��� ݃��W0���A�(����}�}}X����[4Z �����B��z�J	Y0͡�YK�V�6q��x�a�L�;�'�|�#�iӦ9�沷/[mo@P���YU���G����SOu��Ξz�	�X<�@ ?��X�*2-.�1{��xꩧ����o����'!XM�:`�jMLs��sWl���Ou�T�$�"Qe�\u*���Y����x7�nOv��y���lΠ�M�ƨ�O���a�X�+H�:�I�(��"I��?#ylO�ie]�Į�MXi�X�X)IU���sP^b�W1c�N=�D+4�q"�ҵ�W"Y�p?�eO�X��U{_�~�=�̳�[����]���b�>�Q[�����w*F�RP���́%ei-uv�~�ٌ1c��C�t�W�Z����v�j�^WG$��y�˛7~��v�in<����R���1D�H؂���0��lHE��.!�
�s0���"ƪ�U�|�V+o�|EJ8����w�Ց�vC7���B���;�
V3�P��e����aO���Ͳ�_z�^c�KCg-5l$E�Zc����=!ELd1�$ǎ�1��w��E 8=O�l�bZz���Q`����?����Ga)���w��<��D�р3��4`u������e��R�����������&Jt_E4��,y���`��%g�`���Wof%R*�;;UQң�>�Lsy�E|>��Cݠ˸�>���xZU_��3ڇ�� kfbjmK
�(,"�9�Vlm���x����D�2X�a�b�:�k'�Ό�Uڬ��<"U�M�~��@�e?Sk���@�����|5|�+����̣�zÆD�E�*�,�����M-�VJo� @Q�A�j�o�41b��d��Yܰa�G#�C���e��Q�T�:fh���k��|��ۑL��}X�f��A��<]���G�e��M��{#�S���V�N�w�'�.{'#V�sI��Ի�3�e�@^�Zi����?�K8#V���G��GtZ���h���k����Nz+:�=K5!
\�pc���dĮ���r���'��X���O���+�O]a�g�����R�:��M�Q���/�٠�[����
~���^.�εh#��/��PL>j��2%� �����k�Iՠ;ax�|�,އHMl�Kߴ���0�][�Oz��u�&L��R��/�t�n@�����4�ݑW���]Jx�魵�˭�t��k+l���V�:�:�a� C��޸��#*һ�\��f���GͲNFa��_��W�Z���yc.+����D�c=J�G��Τ��x�'����߲�N��m+�����(ø��$!	O%�d���L�)����Xӎ׿���.��~M�{vY�����wH����Y|��^��X�j=���J6�HQ�#�<���},���;,u�B`�i� ��$���m6'+��Y4�VU��� ��J� �DMB������G�����R&sS��t�gP��(7�ئ�Y��a���#7IVE"�-�c	�����'Vo*�T�&��;�Z�:��rs����E^���;���xCfJ�z��bu\3�9E%�ԑ�9�</E�$�H�Kࢻm%��{��=��n.��w���O�'K���*t� 2�,�����2�r��Y���j!6I��S1���Z��C���3;[��
�~yI�b���T ��q�d��	nrt�p�Yȡ�\�gS܇b�&,rM��^�<�ȥR�%T���B���X4�ٿ��6�8���O��R�Ж�;�1٣aM�>��	X[hT �2c�%`-3u����e���re�ɒ ܉!�\k���\ճ��{�$��REf�M�6����9��2��-�3޺e��Z�ܽ�8�6����������:a���'gW����6�+*!3�W�j�«�(���&=h���$��~P�����Ax�22r,�+������c�$��J��w���z�%�lx�Wcs�����Q���r�z;y��K�����|��x}SG�Ut�ܧ^��u��RI�'C���uWk����.������X���Т�T&��~��z��Y��yjgҺ�N�;b���k����R�r���QJ�!��,*�U5)��s V�/���֝�{�]��fd���[o`UT��S ����`�+��^�^Y&>�Չ�Q�ep���l�p({��}(�ܵh8�#Z���f�ƈ*32|y�����y
�b��u.p�oשM��;��$�I}|��u�aR��֡���$�����P���e��D�y�� G���k�7{��h��랉�S�p����pE4K�	}�2:J�7ISNFde���(C�b1��l8 Y�t��D�_k����+S ����,�9kp���:8B+���\勎���+�Մ�4l�pt^�y�96x�]��>�u{�W�����|��=�x���-y׌=R[JJ�W������m&���i��twXx6�H:y�Ξ4�f�3%���L�m�j���tb���
��S�an`Jβ5�l����Pm)'w`����m"t�X=����<R?�&����I��ܣgQk���k�$��!����L���#I)ʍ��ŠeC�i��lLj��C�iKP-c��%��=5�V3^�TR��G����}���;nX�k"	�E1T�о��}�} �!�XUO��v�U�S���ު�5 kp��U{^m1!b�1��~ĺ;���91ۓ.���r�*���H*���>��vj^���Řf�Ř*�m�bFY5�"��?�7NC�=�M�]�&"��z������L��J7�!����&�������՞��ߓ��n�tO���7n#G,�^�/ing2+�VY�҄)�P.��tN#��    IDAT�dӔvmC���Ȱ��/@�BG %'>'0�2�ԑ� ��6�#9WVֹ��P��@K�.3��S�9�M�ؕr�v�N>�J�y�t�UC9Z �e�y2�F䥆�z' )���U*�ݦ'�]\:J&�Jq4�U5�=i��!��wv�\���}�Y�J#(��<q���:s��(�nXu2�k�
ta��C���f'4Ն���`���7n�h�I�gK���X]/���b���*lSmʖm���卖b��� �g3(|��m,��i�� Nlc��j��g��#�/qq�6]���<��m .0(�Yѯ�Yp\T;KՖ��#I%�o��3U�(d�;��G���h�שv1�w����}`�D�hP]*S���T���X�
��*��@z���XwXC*�����VU	PK�>�L��ߢt M��r�6�*pb؂K��zjPu�6E����c;�=0�e 5�JR��er���΃����t"Ehi�X{�D1Ψ��Ř���Z�ڔ��$�^+)O�m����ֽ���;����>��ԯ����n��X���īJ��H�Cb��f�{H�v��ȧ�e-���)� �Da��AR.�n��uJF��Ō�z�Si#�%u���Z&}2s`�k�)a��f�p`����Y%$bu`��TB�_���b|��?��A9.-V"q��}������8D��=��V���@��V����ڭ�,��>7UL^����	&`�0=୴ܠ�K��|ɛV�I��<��jy��6�7>�5�"ϴtc���Mu^km��$�l� )��FT.U�����"a��;a��K�fHJ��������s��:�)a��_޸6VJ�-"^�ǧeb�ɣ��� ď!����_B�m�=��BZ�N�6�{�I��&��|�.�5�ּ�"�kz*X`�Koe�5=b���(�MQl�X��.`E�`U3�]��� 4�Xv��϶���7@����[
����Y�cU�R�T�9��V�ݐ�}���mX�B4����CHQ'��l�	Z��=�I<�F��e�W{:��������ػ3݄�����t��C���8��ퟓ}�{�}mus���j��GY�3�<�������{��-�.�f�
��B
���N���ǡ���H��㭧���_��[�R`U��cr���?���s�Rh�}[�;wϽϖ-]l�y���g%/2%��%N�cE�鉽��s/�����T�V�@$K֍�l��[(���'?�1:!f��/�_��W����{�����3u��n�����7\�pϦ���F�G��Бq����*`U�E�����Z�fk9�B?f;@�Vk6u��  ��L�`3�0���.�>[S��6�]�M�2,N�JV��
�J��ϗeKVm�t�"�5�����n× ��Jg �*q�0.�"Od��w5���`WҠrD$�(�O�%`��U�[+o�稆�Js� ƭ�.�~����AR��ٖ:R:�Ed��������鮼�����������ĥ 4��X{��K^cMR���#�jJ�R�oy)��d�������)
�ڒD�V��ĈOc��U˼��U�&�2EC]}�f�FBث��ߩ�.� �Z�Z1���X�D$�N)�����z��E�ÃZ�F�[�ΘɅ��Z��N?�;��c�7�m/!c8�t�G����O:�z�=k���lTZ_iں%֮��jơ���_�ӽ����(���
��>̾|�m�`xz��|�g�jk������Ir���/�lg6iS�e��`; �h#R����u�fu�1ϲ�\y�-���/_�I�w�H�)���3/ن���W}܎9z:���U�;�[�R&{�l�
��`���T��YE�VZc�6/'|�Y�fS���_��˖-����70�ɸ%�~[VpB凘��f~��D���_kT�p�l�
�D��78a$�w�j�'Fʈ͠O� >᠙6���+�C�ږMm��v
��%�Y�a���K�����m������Ͷ��Ֆl����@3>��58��,D�Poj��W���À�N��r��$]�:+,'xˇ�ݤ�
��$�i��9�'jͧ����sd�T;X"�2/b����3��T��aMj���U�P���@z*X@5�C9�kuoe�5z�ٜ=�n�q��3:���ě�H"���gR�L�X[��s�����e([�kv�t��ܳ�<�� ��8�Y�{�c�(�t�T��4������?���JAL��+�v毜��d��m{	ٱ�#X�o em�z{��g���a?���u��K���3�H*S*����ԿG ܓ5��� ���t��B���"�%`�mָi�]y�e6u�T�sם���/�^Z`����F���T��X���?g5[��w~�d��`b�aGa�����y����@���N?�P��'.����v�Ï[ᰱD���W		]i<J��W�6����?�������e#|_��1���x~P:@(a���@���0�\e�Z]q��.i�A���hӬJ`�;S��>xS�E�Z��S�*`me��
�uڅ��x�"V]�x>��S�HԴ�] !o'���E+������q���`���3ٲi��Y��׬���C%��n�nV�y�+��1�D�p�ƭ��1���D��sG����	jB��(��J��'_��_R�W�uT�J���s��^/�V=*CsY�Μ�����ǘ�>�`�D(	��}W^�A�[��~�*��"�m����X��݆��	�
<c�U�N#��ڇo-�kg��M)@�����~r�j���e`���xgvTsM�s D>Ʋ +e�LC�Di�N�K/����︝,{��v��gZ��!����>6A,$ �NRR�C������-�h>��Io�Q}����C���<�~�?7��щ42�]�Wv �\��T�Tp�>�$m��X�]/ ����}=r۱��e�?�˶`��������k_��0��O~j��٨�������� 돾O���J���Ï����짿��~�i�yv��q��/^f��������Y<��&��lޒ�+��r���g.�}�L����f���%rމl՗\Ir;�*���+pR�N^ڴ�^�{@���V�cy�;����ikؓ=S���ʯ��D;�����:/�x�ޟ|Y�K$�+����9�Y�(@�G��ڭ����61S��N5И>b����O��5 ;�V�Xa7��$���.��������ni��&����}�jꬋו[yK?+��V��O1��'l�'y�=$����a�vk�\�Z��	�E����;�(x��i��"�m��:�ZB�*]ӳ�u�����4`����U��M�����Zu���.��iv�ѳ-� �@@@uJE�RZ�h���\RT�
C� �b������n-�=�"y��u%V�1Ml
}�r�J!��MSİ���G[[I�7)<���{���_�5�3y�	9mU�LZ&��z��'?�����o���6�0��|�+V6j����� �X���Q@�&EĔ���~�����#\Qѻj�L�V	���}|��w�w�-C	-�0\kH%�����k�k�z_���$EZۅZt>���oP
N���J�Y MJ���>�;<��}\�G�a}C����������l�+������\�Y�����iێ�2lB���ګ4M�=>���~�1(��?��N�
�Q�:z�L��.C���6��h�/��I��aJR7��G[��u�����m�74��$ܤL[�r���O��+qL�v`��Z�ڀ�W���n�N�h��D�Ǐ��mn���PLȕ;Jk�-t.����Wy��x�t�y�����[�U��_�g5�j}m���R*R�]�|�;�4�~��:h�Xˡ%Dl\��o ǟ���w�XD�[�5C:��Z@^_�٪;��uhe�9�&ھ]�<��u��W���Ez6�;M��4���5D���X�^���� �<Bl"���n�w�
��1"P�-LvQڰ�}y�9'��G̲�S]p�=����Y�x�����ﭤg̘�c��ɄO�'B�.��Lp�@��O�'1Ѭ�N�������YX
!�������@��Swu՝m�}�*}|M"����Q���	c���<�>x�-Y�����n�����|���j� ���-_z[!EA)��/��JJq
�/%�^T�͖��R�C�h�IY��3A*�Cf�7�RZ�����KXY<3n?�"�����i(=��V�r��q��΢��JP	���=}�(�� ����d��ǫ ���n�R蘏.˳/|���������LZ�����rƄR���F�7yJ�-x����?�[�e%��\G�}'a���vˍw�.6+�R����D�k6l���Z��'.�����jK�o���ü�A�E5�\��WWH�\D�����\$��V���M�8��_w�u^c����KVeK���$�=J�X߉v�.�r9A�A�Z	�V�Hε�Xh<]x;�/���!�fO�j8Y��y��W�Ze��m��V���Q�H�d7j;��2�:����j]s���l�5�!��z�U����J2Q��3��v�I�Wl`���:���O����+Q��&$�İ��=�~����(��� L��X��\蹬)���0��-�n{c�W��q���ԯR�#F���q@(G$���2���}'9�҆�)v7Y�l�$�6od���+�Z;����M�����H��Щ��o�{w]w��|/ihk��9�UDM����>5��=��c�~Ov��y�ƌg'�8ˮ��I�{������D(��f*��1�5��fpl��6��S�8�z��+z⧟|�]����{?�=Fu�5λj����@���X����^�#��3j��Q�����8�J�s`�9�֮V;=R���HǞ}ڱv��Oa�PZ�EVD�Lc$�T6v���w��{ņ*�|�*+ߴ�~��Ϸ/��;r��s�S���m�`{�o�]uŅv�on�{Uc-4��<�^�x!p8���|2ʾ���ٺ�+8����
�R�~6!_��L`���e�-����nqI�d�.��Ga�N���7ߌ,fu,��٩m=I97ӧ��X5ݦ�>��v���n��G庎xl��A�k�j���GX���'������1m�0`�P"`UQ|t����֫�i)��b�*�S4*J��Q��o��R�Q����u����
�c�Xe
ƞ"VG ƞ@��.��[Qe7�1�n��bz7D�b;j1��z��P�	��w���#���`�{���I�=RK�(��-�GN^Fh6�H_���̿]k%hU��2�z��@��ʜ���}-�����H�(q$��p��F]������6ޤ����z���1`R��aO�m���~s�=4����$�R_>����)�NR�E�[���ٱG���5�k�=�b�J��ng�q�o�5�u��|{�	D���sIF���N��$�u��P�1cʂ�A�%-I�8��Թ구�b�w��y�����n�IAj>k��#��u�����K~���X�1e�	��S�W�^w���� A�-�Q�I�-�ٻ�xD��8�����0�68+�D�_��S������q@�3L;^K%ġl�ʿ|�ʫ�~�2
����|����_�B�@��v姮�SN�ls�bw�F#��3N:�>�gد~1מ}q�e�K�RW�� p��D��4��k��������Ĥ�<�%[��I�"rO��n�u�����Rk��߃�[�ƪA�V�Xo���Ǻ;���n3�t e�F�̯yĺ�R�ow����i����[(.�W�1 ���rߓ��R����β�?d�(;pͤ�8f�j��3�p�����#7k ��Tpem�-B,�����jG|�MՑh3��l��i�!M 3���c�@�iCt��	p��s���*9&�ߣA��ۋ�����i�w����{�"�*�l�k���f�D����3%*���iT�j���O?�$Z`Mk��~��Cuب��javh_��P�����ٌQ������_H�T��,݅e��{�7,o�0 d�����?g���"�p�A�9�`��j^j���u5-ty�����y�1\s!Z����@��G�IӚ�Ӛ�g'�Tչ�!P[��H�"&��H[�N��Պ�4�l��?�`{q�D�Mȧ��Lr}A�@���V�#+��׮��直��/�	�<8M��Ն���P�R��-�+Dq�s���J��nL/K�QNGR�Hr�|�}��솛��c�?���Dk�g�n~'2���.���9�t������_��y����䀗��f���BzV/���8>k엿��q�l��po�ql���B"�
"�9���g�~�sWڤI��'�{���|Z4�,dwԇ��d���X	�[�Q5�G�h��>V�X����c���B�_N�&"�3����Fk#��9�'���}��5�K>��9;2�{��X�@�Ʒq�\�SRdmV/q�ս-���6E��p
���3l��ߤ���='��Aey��Z�2���-��h����ڥ:�5�r���o��Ռ���`V�[uT"Vk��Ğ��1�Gd;w�0����n< �D�N>�k�����ttH����X#x'�q�����N�Nו^+�Π��_$��L:N^~>N_k�:{߱�i���6���q 9�1ݫ���?o�_z�K��[VV�*]��K�Z�z��?jC�"k�CQ�v�_�Q�H>�T)��a������b���%-׀l]�tX%��=t����j�d��{�³�Y=��ԅs� ���-D�Bc�D��k4_���V'8��4{�7�5�q�������%v�}�1�zC�Ǳ6E��b7����c��1�&�C�=a��orM�DPD��v���=`u˦l���#��u-#�����߯�}6�G-E(��YǴ����y����$��f2�o䨡���V�$�	�Dj>=�|���S���\E��&j�c��3��e�5b��x��ju"/��L}�˰��,gL�B�M�)gJs����陒���T�L@UӇ^\�(��ʻ�,~�R�Nze-%7I*��.^�0�e�j�O7�=�T�I�m3�W����M��SpZ��-t�0�|��U z��
������X�i�����mYǦ��� ]�_�Gb�*��Z\����i�Ծ��t`�9��fF`���s�E����pD�[�1$ُ?d+�d��&2hf���+��9	���kO�v�X��C4���`}�ZdT�G�Q׻l�������*�ϔ�j�	)I�����+����#��V=�;�Ջ�Y؁�׆��$N�!⡖+dN�N]7�y��'��������D`�_ǘ�N�U�&*����,�5�:욏_l��#ӆx��k',���nE����_@|�{�bO�8�=�XSս�O}�O��g#c����lQsU�j.NN�[Hf��{���Yh�%#�C
7��y�$�&߁۠=[��NU�F;h�L����\m��Ǟ��[�P��fR��8σIk�w�yV����t+�������R�J��Ȳ��mg�v�K:��GD�az��3Y�<�,���^zy��zǟ.�v�\�ů�#����i4{��!d@��=�8g��|;��I�-O�S�94��\��L"V�4o�{��|�^+�Y::B�c�V����kxJ�3|�G��D���"!I��,_JR��V�Z_�E����Y}u�.ዡ-��u�gZ>N]-_2STf	����KҐ)�ȡ�0�W����:�����$'�g(R�4�+�e���+b���#�y79�f�����>��6m8)�8#����ΰGI��s6q#��駟��{ܵ�� q�6�6�S����-)ka�f���N^i�
�6���٨���SV�1l[�$��M�P�T;Z������ x0,�ӎ<���V���h,G�4���|>��^&l̮�-�n�N0No���u��Yxh���,r�?3E&�o�����ւ�t`u�REĻ%Ͷ��}�o�    IDATro`���:S��:|Iٙ��x�G���������t���߷bԢ,��K�\3Q�I��o���<Ϙ��Ϭ=�1c��>[�"�}�����a�Ӧ;K��n��KRt���y�H���k���G|j�ҹ�s-y�|�Y��$dY��7���n��-�%C���̑Nc�B��N<���-iAE�'��|��V�˝w�ݰj]5��3�&�2��}�s/�7[�+��k�U�&P��g+�a���;�ģ�#���j�.����Y�&B��[o���\�A�A>i*�h�ۖ��m�<W?}_9�YE��5�@�/\�^Vhw�1��b䊴�	#�n 1@ο�ضN��q�/Y��P�����N�m��r�e/�zEY����F+�&��T󕐇��U�T���lg)CBʣ}S�ˣ_�Y�4���V�و�����*^6a׳��Y�iI�r}��FD(�h��5 �X�����V�t�im�P��Y�Xe����ϥ�~��G�0���>Ǐ��k��+`U�-�����{*x�X��;�4����[Zs�M���.�����Lj.ꏋ����A�}}h�B4�NU��7�ik�`r���:���a������D�6�!δ�x,Qm��{��7f0Z����PU�L^��x2j=Q�E�I?"�mCɺ�Q��� ���J�$-��d�R.�HU���):o������USS��k����,^�:{F!�={�WĚ��k(��!�h �#�]�ӿ��_��Ժ=�Һw"4\�a�c�l ��3���=�[�: Z��ԉ���ccT6m�lϼ��m�R�E�S&P�!��"��}�Y�R���~�9���:�x�~�2��\r}mܬV��#U�^)����A�!� ���O��і�;�n�4��w��X��9`%#F�_��@# ؎��0r����m���l1 ���ǟ@:�̞F	��Ǟ�M��n�͆B,Z�7I6K�$�5p͗c��X6k�Lm�n�;�����W_N�R7�_�p����p�F�H�����F�Y?\��H?C�g��a/��p�ޱFd^��/�;-�o����F��$�t�8�쭲�.�B�!	��q�����i���mm�u���&~��[��Q��+������!d�E���+�e,eQ��΋�ށ2�Ϣ������^��n�̅�J�#S���(-�6[
s�v@E������R�k앻o ��Wdl8�����خ�5�i>�"l�%̹�$�O*x�3.ڽT�N���ߟSޒw\+�����*�G�M�
�a��ز���9U�Ƞ����Z�M���푝��r��C8ct�7s�e��?i�&�X�W��f�9�.Ao{0u�z�:`���C���ÿ��D	02���.�ZnpsV	Q�&k褾�La��A��J�;��X�"��-}<��UG.�n��+r�G*1��+���?�0�.{�QvԬ)��PM��� �f���,��˩�bX&N�`S'L��f�Z(�JƩ�\gdl��ǯ�VnBp 
L����SI����YQ��@R�%�1z\�nc���؏n��^[��II�X?�)�L)yi����`�Ձ"qk$S��a��aٺ~�}���+? � [�����?�g�R�����BR�\�"8PՕ:5J�϶��b��x�*���`g�|�ע�����$��練m�⥤���:]6�]J������f`��%rH�X(NP4�)���_�+�����cH<�����ӫd!t��p�DFf�
��U޷���'�;k
^���%i�>�[Sn(��5
mW[�%����5�^��O��R�-[Hq#Γ	_F��%![)����n\�����u ,�'���7粜T����ثX�N��*�&M�:-�2�TE�Kb���ۄ}��[Ӥ���w#����c[s��zS֠꣏U
1z���/�R���؜)E�RQkQrK}P_���"JWY�ja������vؙ��ې�q���KQ�A��7���Q���*K����'K"�0���5�h����G���5T׸L���G���Q��k�ǭ�\a�����n���`*B��WS��8n���|��k_�^x͎��n��iB�~2J,�acta�}��g؁�&;��XAF���N� �4CT�r�:���J�o�8~��:��a����"힨�8{��mLݠ��@V#����\���a���c"G����Zg��Roԯ�TȠ! 'և�G������+�08˒�����-6y�h;�����#Q�Y�Җ.]j�v���z�)������ �&Z�A�s좜UM��bV&��������J�-XiO��[��|3|��rکv,}ɫQ�y���.�Ǩ�Z��ԣlG+O���w)k�f��'�=��e�|�+_v����~�׫��.�t.D���[{g�UF�?��I����P�x�"�|�rQ�4�1�R5l��>�GXi�������r�&�����N�@�SF�U���,f6�s�'��3ǥv��~������șwB  ���5D���s`]����T���C����9�x�YC_��X#��Sc�#���n���~�����A^
�>)��_xX)�φtp_^GH"�VjrG������!ĵ5UpY�VV���KtP,ϧ��P��g�5k�7���^�0�V���Jʈ��N�x��X�Jk����#��K��k�T3�C�kC�A�X@ͤ=�RN����66n'��T��eV{�|c��������z�����G0i2"r�t�\�G�p���p�+6YC=���v�1�[6)�v����Hi�b�Z1H�Z�z\�,[�Fh `7q�+ív���p+#X�` �'�䒝�Q� My�t�\j��p��ڛ6Z�j���1QMZ��{��j�ǘ*bm�S�k'����3�8��Y�1�?��YW�1�Ѓ�O8��d�v�wڛ�7�	`��- ;���2�\O����_��0=�ڃ>���k����2hm ��s��l�{���8�~}��b�a�\U�A�ؒ�EpD� d����cA�(��SOt���v��I�7�G}��<9�j�S��`�X%�f�Nߥ�ܦ."H�0��� *�e�"�<��##�<�4/W��U�/���*��h�9|?HM��S~S�ژ��s�Pb�Q~����]��Uz��+�S:>�ψX�EB�<8�V���w\��pR�ٙg��=��P�׹�H��� XcZ�ε�t.Vp}���N�SV�ɼ�+zt)iX+[��XUҖ<���Ǯ^s��t`�����:�G��W"j��1�4N`�UUT�`�p��h$OT�*�B�	���{�,��(���S�A~89�7�x��0Q��X㐈!ƍi��)��H�X{
(hI�i����IA���9�&��V��:����`��QqM�l��2�rK��5�����H<������������MvhҖ꣐��k�^Q��f�E��dSF2Dâ=�W��Lkr��L)�LaZ�n����w2R�sX�����k��Z,�����є��IB&��-�K<��"�]_`BR�3�S�M�"��g�|H�4i$�^'���s0�"�v�A���l/<���{�~��u6�z���F��&�9�λ�/���ߓrԀ����Y�R���'�:t�[�j%�w
r�`oGRo��-�o;���M�g��n���*^�>c���`IWA0�� �O���J�s�wN)��].���{,z�?
T*&[`��D��c�X��,�6�FĦ��P_�h7���&�i�Z��f�C
��7�;�(�@z����pI�F�~���);��5_�y���7-a �Z�/e�rPs��*Jm��'Q9�������*����D�*zr��#�CR��^��;�s���^��+l �䧞z��q�B��Vp,�p~r(�X�������'}`�j�Ayi�����ƚ�}����~��Nhԭ��%��,S�)w���t�ތ�%��g¾T=������Zg1too��K��6u�0;x�i04!+��s���k�>H'��ގ�A���iN�h��� �H�X�������S�WI�N��U��2��1>�|��
k�`|߫C�#8)-^S�A1��������{���ڑ��2�5IFbg�>~���ʍ6�a�'�>=l�6i�p4��h��V�"G{M�,���K5�
ktA	���wb��Ο�42�5�A�?N��C��C������\�f�5�X"ǌ:�"�f@&��$��`�M�$�z�G���{�#�| ���� w�P#&�X*_��i>uGU����z�Dv ���Jވ�g��ѻ4�3�1��s�fPI��C��H4!ʣ�L�2����(�^z�1V}:��e�6� �ɴ5�����AnC+n�E��`UP�`-v���f�VcuV6o��ȖykkR�O}uCJ�}���h��'4��3�8k��]�r#�d����6t ��=����i��J����:�V��N?�^���-d�ML߃�m�N�����{�;����%���g!#㚹�J��X@�4�W{��l����}��Ԭ�!-���S>�|��.i(��QG�ߣ�<Ƶ
?��ИQ�}�y��ڂV�^�X/�`Meז� ���C/��	����0�d�.�M��O����C�gO��T�y���Y�$�=���0����4Φ�� t6gk�G¹肮'%�����hy��G����4jWκ����to����,^]����F�렡oؼ�>C���!�t�k+�	ĭ�T'
P�[tp_[����L_N�{��+��̶Y���TQ������\j����S�R�?C���e쀙�m��3m [�z��~t@��*rmD&O�$yց���S}ߋD)��,���,<z��Ma�;m�"�<����bmZ(1~I��RiBw:�mSҵ��a
-�w��E�}o�"I`ѼD2��T���v$i)-���� �"���f:t()]�&�5��'��HLo`%u3i�:Ɂ't%#���j'@��KN� ��4�R�^�%��J4�!�lw�c�V$��0/Y����$������ކX�n�A:	��Tz�횾ON���d�����mBf�Ǳ�l����[yl���v�.��L{��E���	P�v�c'M�fS���{����3g�M�2־��+p��V�3�B$��aJ�e۵_��ϯ�-��l҃��%<�}|���ͱ�K���MU��x�K�U�`iK�Z�؊d0I�6 +Z��\�R�f1|�:��R�����ܲ��6	����l؈��L����bR�pyP^:�̋��^����[N*�=+�i�SԮI��Yiky���< �#��U�u�	]4f�oR�PS���ZhI�'��R�u4���BkX�q�����mD����q�י���Ci��k���@������������ظ���oނ&��ɢU[m-�-�������~�J]�a��38p1j� ��A*[ڇ����
t�R�j����[b�$E�H5J�`�,R0Y$g��"�d!1\s0����gL�`�Q������O�Y�m%�҉S���'RT��4�`R�ҹ����n9�D��i�y�ͥ�]��k�|K;N$�-���2�T�4�M�	BiEr�Z�[����d�N:gj���܎�ngJ��,[��b�r.RO��:�5Ӕ+�&+*)�ؓj���� ,0�񊼟�X�YJ��r\<S%�g
���Vۆ�MD!�hS�ѱ�U护�n���u���-Z�
��A��^V�6��@���r���+N���f"�!';���G`�^,[�k'm�S��kɣ0����%j�����_�-O�dUa_��Κu "$E6�ŗ�Ϟ�<�+쮻�g6�)D���]����L;®��U��ߞ�����̲�}�j?j�}�����|o7+��S�犏}ԝ����m-}���F�ٗ�"�S0��D���Οw3���<�|��?�4�X�ns뭷"�R�KV����1m_+��^UU�`���o����=��c���疷ر��<2�A�>�T�����Ý*���Q��]�P�)�n��.�Fq�ٌ���� �`�#�x�8.E�a�4>��"wl�f��Iz0!%��,�F(��fN�Q��	Z+p���*�	��%����6l��R�B��8�����ѣ�����	S���.�_�y+��H:q����=qtm:�JE�������:���S��bK����Jā"	�$����m�����OH^�]����5�:�=��=���bwң�5�M&���.�{J� �QZ�o�J�ŗ�Xje�Jq���l�r���R ��hگ���������l�樳�J],�F{�}�৖,E���|�à�8q����s�/�}�#R�ۜ���ʉF
�:ie�}��g�[L�NR��j�����kR51�-^F��{�u�&ҧ�~�I(�W�,�Ik�`־�P�J�M����)JS-�C)w�Z�����见V\� ���5џ�S��A���\M�QQd �rȈ�R���!�I��]����ضa����^��,`a���ڙ�oW|�d���ǉJ&�"ϫ���&`��Z�4�v��^���T���?j�a�McK�]������c��}6{�� �g��g^��o�q�\����&�~��?��PSl���fdW�ϲ����m�/؝��羐�V:�<��
X�!� �-夂����A�bkй�ƽ��+>���s� �L��ywFOG(���0&�"V��K�R�u��ϳ��ZS"�*�$-n���:��$�Q;����L����E���$ߤ&�BSԦ&ҍ�^_�"�kd�Ill�yj{�S���T�u�R: ��!>bH�+���R2���u��M��k[ِ��B� F�0�o��aL�_�7AT,��Z�uW#7��-b�V$�"n�j9��=y�d^[���r�wNOF���@d�P��k"R[��X5q7�2�`�dEe�jfg�a�(��-��VՄC�]�?��|Y'W�豖�;�~��$ ��I��`�W�X��G̹ !-��M K@����JqvH`]گ��2���a�T� #8�y00��ֽg�x���Z@U)aEjL���O�|8%��Y`�LF8oJ�L���K�� ܖ��(s�N	DXsT�'1}�P��gY	_�C�Qwփ���"��L����f����lU9 �A�����RI;�g���K�F�dfLi�~�ۂ��>�;���R�!DM�Ϸ�4�#O?g����K�VB�Q4���`�(����T����>��4�"��w��^r5�)%�ت��S�"i+����T���>f����j/��ѐB��� ���r��E��I'�g����m��K�w����S�(���}>vݚ��Nm,5��
���_��g_�������7��?��i����m�=O����a�|�]uէm�����U53P�,N{�V�G=��n���_��i�o}�{��'�74�c͡�L���f� �?Qc���X�ƍ'����D�nCYbk��Rg=���W^R��"�
�8��,@�GLZR#O�[1� ��������K�]*��I�S7�M&�-��:��7���Ë�
��SF�� �3�c��1W����^E���E+ચ��5
�
x]�p��"6v�@��cl��"���[9��6m�6�FzF+I��ɕ���2dL�3 'aWF����7�Kr+�e�?:�5���_�����u�s����&[Qو5K��j�C�z������*�����}Xwuwv��ےRv��5Y��}��fC���"������v������k)J������tT?M�Q	,�xt��I)]�tC^$q��|�[�>��]�< �>���UY �+y���K�S�ȃ�m��f�)��/<��JۜҢ�ꐳ������窈�~��9�����`�e_���GCn�L"7fCflg�a�O����GY����U�֚�fm��NR��ѷ��M�[� ��NR��лwEϚjp\vg�m��� \�` ��g�b��t@���`ަ�����mˠs!vy    IDAT�{����X��A#���A���������
LH�����>|�+����5�a�d�ev�.���P�"-?jx�=���vӭ�3�o�}盟����)���[m��}��߸ڞz�%{�������ȣ��\!�A����Oѯ<���?du8��$l�@���P%|���1A�F�H�*;�U��f4���_�t��z�cp��ƍ9ʖ,Yl����}l���z���B��}����<VM�iހ(`�Cy���>����5+ ��J�xZE�{��|.���Y����n*�(�ż@�z���
L�F�4�N�Uޘ����[�`;���[��q�(F#9 ��Y2L|��&Y�B�o��H���i�w\D�&��x�A���3��5�t���99�5S�����r���ҿk�дi��s��:�1%#ڸic�Wm�Ÿ��T��j㚛��P˫�PI/5��� �I���ӿ���6T�"�=[��8^Nd
�$���;s:l�d��c"HP/�{����UL���꽁UĒn�"Cr�0����s|6�+%��L�tr�|���Wxv$�-� �NdIv�v��B��`�:\u8���0`#�,�TD� Q��?+����)�ȡ��`�3e���8�t�nA���M��$@�"�U��ݯo�gkZ�YQ�\E4j�k���X�pi6;�9�.�ڙ����Ҁs�W�3;hk!��y���)�o�yL붜B�, ����5��p�T�~6��ռ�J��³l��C��V�|�~�Y�flG������Av���ؽ�0�x�;Z��T]�U�P�?���'���@�"��m��`�6��/}�~��w7���x�d@>���4�H"�Oڼ{^��CH�5k_��.�?�z�=���]�N=�T��O����f�X���h yv�5���:�����K<�� ͂r;��/�[n{��{�	JCp�ⱝ�l�秐TQK�J[0�V�a� �2��Kc���7�p�^�[У���mM\uVE�V��Ucm��T2~��<�����S�X�2U;uƬ41JyPy���O=x���x��L�*^��~T�&����3��|�7y���Zf�X
ۀ��RB�+�M�TjQhGv̧_8XM�,d�r��5�G�����`i��Ҍ`�z�4�N����"6UPI��G�WХ����"a/����S{��`u��H`Dτ�߈�\A����I7A�H�2!E�,"���p*c�"�����WWݓm�C��+���Pn�N�N�)��=�P'PtрdR�����b�^Wh���O���y�;?���$�aE2W���.���p]_:�)�Ԟ����=�{x^�p�#y/:�=ȉ���}����=�J�p�)pT�w�@�<��D1�6ִ����V6���t�-E2���3�k�U9m�Z�֎<����S-�^�z(Uהn�2r*����E����~�4!%���6�;�!P���k�Pw[�-N���e�{��ʆ��[��>��s�)#��,[N���T+�ũ�䘶�R{��E6��Q8H!Gp�v�;�n*�i-�D�#�ɤϔ2�G:��� P�#{Ld2���}P�d�?�����׾�O�ڭ����� �!N���'.�#f���;�wﳴ��N����LC�w���VUO�L9��q>�gφ�r���Xg���_����!�K�T:s�f9�.iH��6�� 9�y����Uc��x�.V�� �X��L���%����mf�v����c��2��D_tME�����ў~�n�[�
�+e��2�\1Hv��6�~�n�� ���F��$$]Δ�Iu~���l�l�F"V��$�4��q�D������~u�+i�Z'�M�a�Xt�p�v!�aL-��l��!6}���C�Ȕ����Y��"��&��S$�8�/=��T׮z�~�/P?=����!����m�D7���k a�(B%'̊�S�����	L��J1�4'�9���&������Ťu��7�rO���B�����І�{��H������nW��_5�ß�s�}��%H"W�wn"H�ɻQ������p��#�£��ҝ�����A���f�H0e�l���6y@�͞<�
�@�qb�: (�d��ɿI�������͍�tc%�E��4�#���k �����C�o[�͞>֎�=���K�U'e�
�2�.j%%�О���u��d �)��t`��2�[������6�G����T�겳O�æ������| ,e�d; l���yϼds��o�L1b`����cw�Kځ�.Ίd.5d"�jٽ!�%L:�;d�m���s3e����3�]����ؽ�=m������?h����B��$��kW�0�$�cv�y>��S���u�H{e��T�F�YP��(�%�b�cr�aIA�@��9�=#a�Ti��ށ���,����KW~�N^z��믿�[�߼��UY�iS�q`C\�`��۫���)kaf;i��$5�/R�>���<v�խyՍ,;��3��j\�R�R�P��Eùi�q�Tw������ )�v��Z�iVc�2�J6����n��^C�Hx]�i���NZ����ت�
�U��c0�����6z`��2��Pdi�b����C�Q'K��L��:�nh=Ft��|E!J����Z$���b���0��8����D�,�a�,	��(����3pūd �G,���I�a�QN� ��ʫe4�ѫɾ+%3ii�j���\������>����$������Ap��s��b�&�R9T��$��y�0,����1 L�P�Ӟ	�"\O�'�4
t�� !\�[]JH֨����v�z�N%Zʜ�jH���c�*h
���I}du�r�Ľϼnw>���l��9�\�����2��:����9�p?��v� ��fzH�Mu�L�t�^�WIX]�b������:jM��L�QqtÚ's�}�����R���\ߩ�����3@�d��fȢ��\lE���l!_don���4����-�-�mN:����i];:�*e��#��I\mz��u[��6j�;h��m0f����z���oH؆Y�0%C{����"t�kj(�ᰐ�)P�&�#N�t���m���)�l����	�\I9������0:�X@_�P벝r~D�)T�u��"���
^�}�崵$����W�XfO<�sqbq<�X�,d����E��\��:۸~��,[��N	D��l��X�	ŧ}�y��ǵx�U�jB�H(�cJ����r{�V��U�����˽.����3�c���Q�Q�v�3�%hC{M0��p���)��*�[+f��u���F=E�30�4.H�+ NC)�v�O/K���(�56�!�Զ�̛�$`�u"�U��3����`VR��JT``�ih��G$�u�{�=k��4(U��er��;�Y�J���c#^7�(�D�8
�:$J�����"6��b6k���7�)���ㄇIQ��ў*^��<_��uN��"�$ ��"=�ە���1������h��=�5�
8^k���D�ǲI��V߫+�(C��%m[�$'S?����HQ
����^�lE� SU�X#�껺����&�]���W���w�r[�a_���飬��b�Ze�����G��ϖT���Hf����?����X�;��=:6��A���L=Ȯ��"�0b ��*��g�[�b<qL��o�[����#�n����m�Q�`����ֽ��R�qg��O��0�+�#�b8|��8��_��mJ��t,��Xv@��V�/���)�58)����{�������g"�%���"Z���O���:����`�Ȟ�i���==-��_@*Zሂ�溪0�U�p�dQ�."�M!���=�x�X��p`�j�ż砍`I�u3a:S&ק^�N0A���P	PNP��M��<��,�w#���>q��cUJX��}����,�����8��Ƚ���ڤT��m4�\�b��X�j��ޏ���2P��Q���K��c�K���]r�%v�QG٪+�]���rOպ �S�n<ՉF�Î����Uii�G�K�HW�X�g]D�:�j9,	�#n�X#�t���>����}�Q�{r#U;�'�~+�D�_�����'�Q���#:���՚|P2�/��U"��X��A�e��D��.l��5$Y�ભ֑�hƒf��U�![*�cxy��@4X�'
;��#o��4��nՎ�
�J�#�]*r�9�I�Ǟ(^�B�;�|�?�G��=�*Y71?�3��ה�'m���Ep��\9\ZA���Lw�I��B�y:�����.&�OHw��]�6����_�u|�mK&�#�v���ὺ��7��4(��oO*8���lOlų�j�80�>���� Sґ�##�s��f����>�͚�,��'m��/R��� P�wrt��RK�m���#����>@+Ғt8��~��&��p��N:璚mY��g�?�*��aoX�˥ev��Q���$󕩾L�D.8����#i��4e��A��1<_�E�@� ��Ek�o�k�gԊ��y�9����A�0_�>�W�E5}M}Y��t)���^�X�=ٻL�GHz$Ο���%:m*M�QsN�l���$ߩDLl����c`�I?�kk�n��<+ç�Q���M0�ɗ��2A�D�-TP���F��s�5�f2���#��(&j��2��
W4ѯ aw'��%�,�.�s7�w��N)_���kƠ�Ǫ�G��]�D%��v촏U�z*kys�qt��XC/=���|�W�?2� V����K>�dM���l3�01�S>q��N�4�F�	�J�ÍT��g}��u��&�5FR#�Y����o�h��ꑆ�+�U�Y?c���\�I	�C����������|����V1�hU�!R�@u�<�a-�H$��Y�T�j}w��čۓ&�xG�sW��ѷ䧀AT�V<w�1���D����{
;3ﶿŽ��ʎ).�xi��TOD�A�j�Һ�Jϖ2�Rbx��^��LbО����v�?�'=%鄼��]�:yp�]u���$�ڑ�l�:�X��4�x�J�v�D,� �09����9{b �*�_�HU�����]�o�l� ����<��,Mlq1�� ��aLUga�˺6�Mw�o�>����O�R��-������Xԋ��5KQ Q�'
���j���2��K5J�T�:Ɩ���d\�ïn�_��W[[�����ޒ"qw¥��(/Yge�D������dR�,!=�~�GQ���ܿ#�˼"\>����t�8�	�5=��r!�����s���gQ_x�!`�s�&����D�`���F�U�&b���`=-�A�يV�&�]�X�vn��Bι�Xܛ�������{o"��ʽ�iIƽ�>�?t�y䑶�4�����|��MD�X��2e�6j/ kOV���!�?�s�	)�KRa�U:�*2M�'�zPY�c�����X=R�|i�z�[K�ǘWC)I}���{�_wR�o��8xj��+��HYA��5�~��5'pHX�1�e���㾲����O���î���3�!�����F��k��噓�k��� ���* u�(��z+���};'{�^��}v����ʱ�^�~;~�8�}5�P��q��oVbE����W	X�{`}��V���X��>�����h��h��9_$}\�1F3a���É��/�R�]"�,JQ;֘�����8bE��y'b��y��q� ��Ji��I4��nFE�ޥ��#�m�_�~��E(#O�Y�&�I$L���]�Y�.�>��xyn�$5�P���V-޷/���&��L�B�zw3�d ����s��.!hio�t�)�����D5Ω�ˑ� �(�vq ��k��І�L���ng�%<]�]�C��4���V�"V8�#V9�X�[�5�~w��1��6i �f��U��X1b�E�0�;�98���΁��0�l�6('%@�`E�Y�K�D�	DZO]�"c�.%uL$�1a���oz�,2����5��_��&����rx$k����O����Ҡ�̺���&�O�@�>6�;�k�]W_�^?_����}zV�{����4�?�d��4�]o 0՚02�%�mk�!q|+x][Q�sLXC�=P�ǭۭ��XG�d�g?�;a�X�nD�:#*�H��#��d�2�:+������{��~�9�GN�Q�i�2E	��
�	�~��m�Xz!�,�J��\o\���x��_��i��;���ڞGm��k`�h5v5t�r�e�� ;V
�8�5v�I���8`mGY<�PI���C���#!;a#�a=�h����uS5y3��*�������6�T ���""˒�� KZ�^wO{��F��zgWp�*TD�޵Ùm�B嫢:&���ʣ���7R�)�����pJ )iй�D���[�Ju�{~�9�;���qT�*"�f
{�:�F������#v[ce#�κ��q>�Νّ ��DZk6Z��X�-�������>�4����w��!�*��
X{o$ݔ�K��S�ڰ�������]�4J�g�&�@��b����R����:^�O�X�W����.m��F`��I!�R�<�&̐N
p�!V�Ǝ��$��Y��)H����uXEB�F��ɑ	�E����������Ġ=}��iS��l�Ѫג`�*�ҼL�)F-��N�zUE�"�)bUk������uO�W_��3`�V��ࣧ����j���)U�#�H{��HZ>��F����ǟ��h�H�I~��Q�h�4U���/=����y�I���TE���ʘj�d�^�����| K��O��XC�������8b�O��$b=�>v���`UF�т���p�q��8��>��Z�2��5�Z�p� )j��w��[�L���jOQj�}X٧<Q~��G��3�~v�\�
X�Z*Ð������bʎ:����� 2�<�fWy�v2e/�{�@�I��&�m��8m��^�K�6�u�_oq`�<փ9 ��*g�v�^L��j�]YT%��<��s5����*3�"�����X�o9�^��{ �-Ll�]t�]U�O��z�ތX]}%-]?�[�8 d�w��
���"$q�|#󐷧�7W:�z��7d�P����r����_R�Iհ�%�jNZ���eV.�jZ�4@@ /�&EЪJϏ��TlR�da�T�� ކ��(ӝ��&����������"��y"���M�o�\��a-4ױ��u��}�p�x�kW��bx�Z*�gJ��=`����Y�ulI�]��s��}ƒ
f����X�"��n���2�U�D��<aw�
΀�ڢ�6�52��d��Te3Ps����X����Ő��dCD`͠Ģ������m�f!��WMU�ӝ����Q�����Xi��o���egm��fh��$]��#j%|�J?AĪ�*JDE�
i���4�=��&�Y'Mw"�<N���#8!��o�C"�e���>D(s�۩T���x͵UC��b��"0�6�,%u7��Ah�էդa8^�����C 71�5mhW�.��s ��{�/���}�D�FqIR�Rk-�4��KB
~�5FG(�T]WZri�92�cU��K�
�65��"֝ ���x�f��i_��=[ /�1���uG�x�b�!�҈�c��&��ٔId����p��Wo/�������b^v�������{% ,����e�S�1Z���X�y)����ˬj�B��rt��r�w�ˆ-�C���T#RY,���
p�y��n �� 4�Yn�up�X��.}��Ĵ�u_}���C���I���i�mB��J��i�p��Z䥾�^�����
�X�)�O+bu`�����t�w�DB˛�E^��^j��=�}��V�TG��s��2��l��R���>h3Ɣ1���U=��;���.%����Ӯ���
n�ƪa J�a�X�S9���搕*�{z���c}b�Z�B�O�6b����"�T�Q
L�/Z+x��kn�޲) �|)��Tc�G�@�C���T8���b��    IDAT�h��f��V���c�= �*���=��$3�B:$!t0�A��)**z��׋z?�EA�	RCi�'�齗�Lf2��k��̼	I&�ϗ�ޘ0���g���k��=�^䖮^f?��G����t���9��z��[�ښ�F�B3���)'�3����U����i�M��=���3�����5[�6������稜�A����������)��/8`�Ƞs�=Jz�Y��:>���@6&�#Ɵim�%�>�n/c`�Xg�"�h3�#��#Z�[{t�h����z`�8,����h��{nI u�Gb�o�&���ޑ0���5ʷ|�m\<��e�0����$�r 8@ǿ����}���$ʉ��p�����%����ߝe�����&T���Gc�Xs�,6
՘�Qp����|2V���/`T�Vp��I;��g{�P��շ���>J,I�A]s�<�G��viC;��\{���֚	�Y�u��?'�soM%c�U��3Vѽ,`H��^s��L�*��`�\ B��#Ņ�(�w�����z�Q����ݡ?����GEl����Xi���'��q���c%'&��]���>�Mο��9�����6���`�J�MFv>
�(~9�%:��O�,�ɞz�9z�5��<S)g�����\��6�	h:�:�sd�������G�]�;�����Q�>g��t)q�h3�'����Oo�;g&��P�}N:n���k���7c�]��=�G��*8 �'�J�%NPEv���1�|�͚����/� �f��?�F�V�+X�K�
�1k��2�
�D����ɣ�2���W��څ�Q}���]`�r��X�����?�oo��hT�u�c7#�<��h��ֻ� oD^�l)gfN�́��d�j����x|���m��B�s��{�����{V��~����;�36W �"����7��@ukJ�|۴b��[%2�'�uD��B,#s��Us sգ�,:�Ω���L;{�]���}#��!D��ܰP�r�r��m2�Ѝ�2��eh���Zknw�lɴ46�V�~]� �T�Ub���z��r���N�@*���d Y��d<}�{K�Jrp���J��ZI��5�м1}��^�hk�MQ`)���z*�YL_�B�ᓎ9ĺe�YςtK���#��=I�����#�[Y^o��[a���07w^���e������c����=$�(��Oc}N8� ;{��� $PL!����j�H��"�[�zoJn7����n����0b��q;-���c>�������?�q�*�±���!�]���{�� �{�}d��.�dCa#���b��e#F���+`]°�$��fpT�m!������HP�GϞp�}��	��'�3/�j9�݄��
��\>�n.�!��i�܋M�Z�֭�.��k>6N^��nSIm71�����{�����+8������V��kl�:��K;G��p<̨�0��f���� ���m�5�o�F��e˖��O?�`=��Sv~���姫�u���]?���]�rvV���u���O�̞C��a0��>V�!3�N#�������B�Gx�*��U����o⾙;E�y:�(�	�����.�l���r�G�s�ȂZIf��ٿi@@�b��S�f}�R<���]�~B�mv���+�?h���>�BA�2�\�=�=K����ٶ�9���������3MN��NBMnI�`t*X�}�3Mgǲ��{�xH�JK��n�v�٧Za���J�$����rJ���fw<��ͣ�#%�lF�q̂9�,�e��C�J˦�v������F�,op@G�-�2���Z��K*�l�F{�me�Y�d#n��C��[;s�����j���X<��Y�Q��
[�����9��z撵��R[Wۊ�=�7�Ј��=� ��/n��ux�V٭��A�Y��j�ۓ��bb��	!�7��C����m\�ľr�v��ΰ[n�h�gΧ	�`Ww$��J䢉d�ݏ�!�<��b2��3ϺO|߭M�j���ICX�k#`]jӞU�:!���ܹ�ہ50�]� �Ç��ʄ_��m�*�8載�%M%:/l�n�u`=�;�~fCm�k�aA(s�AD:^����g��:z�h�+):Peb��E�������n6y���c�¥�o�Ӧ2��.}�ΰ��}� "D�;��;ب��bb��<o>����w�Є������A6:���+C�PQza*"%��l	�*e#�'i'3�KI�cץ�U������cس��νۮ�˝}J"á5�u��~'�sCfc�V��h�Md�y}GP�R�iB�(ʍG��u���Ȅ��ks����g@A�' �lx�t��S}ģ�G3|%C�P_�;�e�:ԭx�i[ZM�q>�MB�0;����fr�4Ӻv�ؑv��_ #,�٧$�n>�@��Z�E%�x����Ǭ�qrSf��-��4]+�ץ,�ٌu����5c!X�Xj_�p�6b_k�(�2�w)�hO�n����J쑗�懖�kԪG)�ݮQ48�`k]���k��{��?�I��Y�{�r����UB���1���k����}%AR���k+���.8�~|�=�т���T�����DCR_Y�,���S�������=�����;�Y�j�Iu k+�B�y�D����=hmV�Fe����kt^��� ��^�,uG;��U%9e�a����OXg���[f@�\��KLm3j<VF�_w'�K1zW��5���|��d{���l���Xۘ�
�&B�E��Y�v����;���l�6S%mX��h�[e������&�Vω-�����s�# �D�i�ٔ
�q�,&���L�i��6���!@��\��6���V��P=X*-}���Y��#7��*T���@M**)�0�K�0}�T{w����	I-@����t�kuI`MC��}�+��% +�lw����w������R���7��q�,��\��,��V)0���i�ciƜh+�:��mqM��a7�Fp�X
L��9�G�`�a�I��� 2�Ngmxg�l�4.���G)��P����V�8�69��c��7� - �~&���P��w#DL�o
�j7ZϔZ��cl4�Γ1nhP���둢�qj��Y�s�?�G_��L&�5X�܍��T���x�o_ Q�k
���U�*�$���*�Q���ե��ﺌ�8GM�nw�p��7N���գ6#���fșb�P��c!��qGiGu�=��?��7�a&Ki�##�A+�u
\T._�q�22������o#��1`��f��Q��:��YN���5��٭�^��r^��*xkkP�},cXS0�.)�
��͍��E	,j��N�P��Ŕ�n�a ]c�֬���1�����=cMF��6,�a.1g�|;�(F���
�O�GL�vd1:���G>�AW�Y����ls@m��j�Lļ$ԿZ��Yx��Z$�߸�j��M������ͷ�s(VS�_����o���I�������U��v�)�x��Dm��ߴ<�8�6l.]�X��5T+�7�'�
�������e�!��Ҟ?7{߱�3 �o#��d���K)#�j�T�l��#��ƚ�0�5dhxp�-� ���(E�?�k����@�g��HT��C���O9Β��X��G�z�^F�\S(��������E$s�'_q�?�3����vO����R�Z69��@��Ib� ��E4k��P�j�E�+3����́�΋�pY>l�W�;���m�X�����o���`���`ݲϡ���3�*G%�(��M�RQ�$��V��'f\x������G�VX:����^䏦%���Т�1te�V[	c��p�M6y�:��mwX:f/b�Úf�{�*`]�Ħ=:|��|�ƺ5*8�裭���uˌU��3T�Nk��*)�ࢂ=c�?�EƉ��5��Ǡ�TC���Dխ�d\w�~No��l:�r���a���J��kP�m�+x˼ik�K"��Emz��؜���Rs�k������(�ݲƺu`�@5:�K�ظā�����]��ׯ��J0�Nb\Ӭ�3��w�uz\�h>j����	���߉�ygk��������i�84g��:����_:ѿo
�}�-{���-93��<h�����T���%�	�� �.�6�����o�{�ʹ���og�?ƺ#���UM;uc$��E7�B5�
)��-*c�#���W����t;��:����p5f�����,	j2�l�_C��0�VGWnQ15�J��}� �hr��_#�eHVڂԳ���m�-/���*�Nݴڮ��+>������6eD����  /�Fzk��4ٞ}{c8J��R_*#�|��*`5�u�x)����B��2�D`U[`��v�zFl��d�WU��I)G�1Ԋ'�?�N�0��p������|z��N���x{�-_���%U�ϔ������|ڑ���^�קLua���e���8H�R`"r� �$^z����t3`U�����a�R2�˖5֝/�4�a@0��~8�Y����
&V��K#�u����Ϗ��H���5�mY����L��Wc���48o��2>���D�X��;1z��kG��b"�E����R�����a6��U���i�ia�QRl_��������[<��E�!7��G��(_�U`۝�%ގ�Sc�,	I���=m�*S+B�^�m��'8M��˷�~�~��${���3��0�,ه3�ړ5�����?O�Z�;��#
�3��5�]�Yw�uN�J�IR�Y{	�H3e�A����SW΍Z Z�*�j���e"А����ZudFڈf�EF��o`\܈}��Q����J��v���V�"�h���Lוe����?�2B36��q�&!e�y��CSt���vX�^2�O,��X�K;j�޸�@a�n�Z0٠2�6��4��T=��6u^��817V�%^X��t��׺&A���xIӲZ�(c�3�����{�E���fp��=�P;|�0�U�d={dڬ����{��ؓ�>��J�/�a�1�I` k��|�Y�j�?�g?����m��2��3�ʱ7�]
A�T��XX���*807��2#)��:x�S�r���1�ƪ�q2��#T�����[8����%ȑj�Ů�5��_V2���}��@$���h`��}�D�>��&��.L��R����
�ب�'Xf���U�Qߡ P7O|���7]�~҂�L�MR7X0��#���.���dxM����=@�����=���o�-��0��1�cf�:�3+R�E��S����Ck�*���Q�]�MF��S�h���f٫�&�'�x��
������w�
��I�.��gfR3�ׯ��x�Q=������p`�n˲|T����iwQ���J��(b=d��X;?���3�AX��UX�5i��Mnt�\	��܄��zJYZo�tY�q��$�SM5
2��8V��j��5KI ����x�@�� ;��L1n��F�-��-Эx֦�������;uEz)+|�CPw�Ǫ�H���Ҟ\���H�=�G�;�;���h93����I��Y&V�nb��r���D�*�+��H��A��6��X�Τ��SB'���J�s�;�X}^�Ǻf����c=�Um�,�����d�[Sʘ7ܣt.�����UWٺ�+m���h�h+�g(���`��}`�֓��py���۩�J�ؙWp���ox;��A���Q�X�+?��qU/����5U��מ���
6�袋<��:j�G ����'�]P+�5Y�5Zhs�-�t�Lƚ�G�/*h����a��۴�<F'Ѧ�h��d������&�p) �n�6
��h���6��.4|o*c��&7��Pu�Bg3*N�d�;5�A�&��0�^7(�č.x��޲p�HE8����?���6��K#�k����)�oDC
E�o��ÓZ
4s�lf� �d��fRwZ�T��v�U�Pk����#����;�&q
u/&��ܹ�_�١��҂�a���m����D,���|<��޳��-Ê�ƈ��J�/矻ܿ��ۼ��CPGұ��3���#tpRU�@{�/��Gt�F��r�݈)��"�Z��qj���y��G���6�Ye��Q"��&���1 Q=�~��a�"C��'=����;�r�ڋ>2�1FIt�>2�؋�����Q��������Y8��Y�� h����\�Ot7����ک�?�~����r2�%�c1wu��9HxH>���B��M�[5�Mf�&���8Y����,�P���y�g��l�����Η���y{�Q��JS��ayW�b�wW���Ka��[YY�-]�PJ<4�����Z����=՝�A�֬��Y���Y�_L��#k V5ag�
T������X� �+���=g�MM�6�[n�����o=B��2Y�N��Ҧk�������"� ��5���~=�m��D�n�H�-�^���X�&(�ToXcC{���N�Ī�����ޛ>�V��D�W�RC)_���e�@L���Ӎ"S��VҤ��5oI��3��kA����T{yj�`\��{�!tX���V��Vd�����'��v9���`�e.XhM�����e)�{��!�������:BT�]��ʖBӂУ��]v�Hɋ����<�^}�M"T]��ɘ<rf��>�Y��9��e*"`�C�w�{��K)964�9��B�T��Pl���╣�2�`�y�����d͟������J�Ҵ46����7zx�+��CoxD%��2O ��΂���C�d�1p��E��o��i��`����P �&�V�R� kr�2�HfA"�&a�� +�o��H{Xu�[D
���hwifR�ٷa-��6��$�a��9%�I)�Ǹ��	g�ϋP(���(ٕ0��`}�n�ߋ�7��̺��(��Ev�����
��Z�m]�Z��텗_��*���ڰ���}*xW���sα��:����^�jU�M��D;ð9j�ԉ�^\B�Qo?�r�b;��3�X�%{��+���p�Q6|p=�f�箲��|ǖB�#�:��cP�nU��+�y��>��z�^}}��0������=��V���#�)MDV���L|ڦ�Y����_}ť6f��d�&wf�lQ������L{�'��a��K����e��4e^7&֗V��|Ё�>oϒ����T�¯�)@��2�9�&��i���+����T2`/��xǁU��)���9~�<E9��w�ޮ
#�H�ͷ&9�fBu�C������oNx�q����٭���aK�%�6'X��zl^�����m�[�/"����&��0q#{ ώ@ �J�,� V%_����^Q0��d"9��Y��-I	���Vؿf�U����Us AM�ly��`�Ux-Ǩ�O9��n�:�Ň�U^�6�_���ѺC����_tFkѾ.�(�U�V�{L��
�w� b��]�s�=׎��h���v뭷��������p��E�~�;�:��~o�Wb�%^*��k�2��DF:|@"�+m��%��>`�<5�>��e�^x�����'Z�Ƽ^�(FO9�x;���{_�g�~��P}����sO�	��6e�t�n3_ˋ/��֗o���z�U�[�E����<f��|�̀e2.Qy�1���iLɵ�u�mĀ^����
{�i��C[A�ς�%��ג�+�֔e����`�3aEsZ@ k."��d� k*�@ע<�UpaAԌ��o���G��9Rb�i}�����bC�g�yfD��6>�:�༧��Z������ظ��"��(no��y^!{��mNm�wߜ��h��˺�q��T����d�
�Dtb����-�/~���p.Fj��0c���ȍ;���&�lmc޵@2eS�w�x5��3Vf�j&n�y��{�6E],SdL>`�ه�+c��;x�Z� .@-P����)2~����۸�}Қʣco�Q�;ei�ǁ���γ�:ȁ�O����몉���I'Q���=k�&9G����;T�ϰ�j�d�.v�l����A��Š�n�(��*��]c5��7�
���qa���P#�8�����J�b��孶b�*��'�g�`����3ma'���    IDAT��C�j"��o����Sb���?X��ݸ�?����G����_Q�%#*rz{�6��:��C�����R�ǣ/�C�<f�жu���+�*������R��&E�qd�@���Qc��A�5V��e���P����T��X����dɔZ�]��GX?Z#�ل>Vm��^���%�T����p�(�fܓ�5Y5֠��K���6��f�o����v��-2�H_���1򳄩Z.-�L��u`N����W"��JC|�OD܊������>Q (�Ϛ
�D!tZB�Y|`M��<�ےpGC�-�$�`<���F�![X�gǈ�0���I՝\��Xjq�;l*[a3�~�қ*٧�4��M�*�i��Μ��݉B�:�d|�5���?�;���UY�A%�fX a��Di�M�=�Yd��yV���O�:��3�{��j��d��m��� �y����kMi�6l��?7�m/=�������^ kzDCc>݂��ӏ�s�o?��=�<�k�3��N���~���l�{��e�\u	�,���'Ȅ�Ė��G�(�i��R�Ȱ�:��g�/�=�^~�E3��������M�g�SR�բ����;|�����"nT^����Y0\C_�(!��LY7�3V�7h�`&Vdy�U���M�D���L�~�����X�F.,,���LHJ7���K���PWM����-�a窱�zc�����������PQ-u*V�ƻ��-|�}��q�Ds+Yj{ WBQgA ��]'eR����qW�g���+�����@|��,4U"%u%�*'=����*L�r�%�uj<V?�׸y�΋�Z�=HT��Ӽo���4< ��g�nm�]�T�%Ϫ�F΂e��	�:/� �	�Z���Ջ����yI��w��&���~���꼴+T�j���Uc��)
6l����J8��X{����l�1���6���X��"�=+!c�����e��حw�mI96t�`�ɍg���jO<��'��*81E��*�C���:�0;�L��[�I��L�����N����[m=�^�О��쵗�سϽ��x�uXr����k�v������A�K0�ƞ�KV��ys����7\�d��2}&2��lVt��MAi��wD5�9v�	�_[�kB�.X'k�P�%��7 �QD�b2u԰�(�4�#�A̟�K���T�Sz��`U�F�WT�&�]f�!�ֵ���ɋg/�~�W��}�PGu��J�c$j
���#�o�"?�>����|5\�{�U!������{�?�ݶ$���g�jk���Pɱa���62S}�h&��=FL[
{�wG�&9:��Ч�C:�X�fe��g���M�l�:w��8�����Tň��ڌ��|�%��묒U�e�=ULf5��i%�m�)��>�~���>��!	�W��u��v�������"rH�����㌵G�^Y̙;�*d�O�zTp:M��Уr&i�*��������͞��n�����;����]isf-����+�/���l�˳����ʯ�j_8z�����m����s�D�z��yϋ�
e�؃��q��'y�&B)&e�sA��[�o]��g���mj�����Z����=��+6�	�p�e����Ï=IN|/���@ ���sS�)ݸQ��k��SkJ��-��v�g����49GT�v �UYGv��GT� ��2>��^��@��&)����r<���i9��6����U��|_�%x�կ&cP��+��-(zC���#<'4EYg��hݜjb�D�T��VT����������F^�ѐs�Ec�s�\ܳX(Y�T�$Oi��Z,�nUk��CZ�-�kO4�@���a���h�ڒ2I.�6��i���w�{��X�}�m�umܾY�nXC�(t�V����Z6�׎N�鱽�uk�*����dd�2�Hl��dڍ�Xǌ�Y�_����/�H�&Z�LV�^Vҽ���K�,b�542����D(C��L�����̊����y�͛;����n���=��ҳ퀑�ο�d����EY�kF#�YD1���B���}�6�_����3N����-��.��M���q����ٔ)s�/�t��	�]s�?��ϭ
#��U+9�����;�oj�_�瞟l<��[�i�D+�ZZ�߮��{������V�N�����X7,�ayj��dJD]�������k�R�O �ݬ��t{���6��6��ݜ�U���:M�#�be�Z��i�/�o���L�`��T�Ie���
X{�mv�Z|�맳l-��s=��Y�]?���t�tC����,4�<cAM{��Cىb5�hлW:�t�1Q�z���ow�RW���mP ��2����=��Nn��Az���3f�~��o���~�6����!R#m�#M�i�MI���[$#��s)@]ċ[�(�`�w�^ݽEI���J�626&1���4����,1�Y��L%P�� +�m4�U^��h�����qb�dD�=`��}�X~!T2{�G`��N��i`�9~'`����V;�}7��xI�ΕE�y�.
}�A-���8�K_T���K}��h�|N(f/�=a���j�GK�^��e�0�����nU�=��6{�jJ���j��
����^��+�ya|`סv�Qc�~m���K�Z��N>+�S즟�c��,��\����/w������Yk����Jjw?��A�fۓϼjU*P���P�-Y��M1F����Ưً�̱�����9��z�"w(�hŷ��"�#���м�<��J�;���O-A�Wz�*yyyN7� ���K���v��m	�;������s��C7�Z��$h�eI��ƐsQ���`��hH�^`��,v��l�m��:$��������
\�4л2+���#q�L~��#�������U�x�i)4W6�Ɣ���g8:ɝ.A�� � �Y�� |B��ng���@���1�vĘ�툃����M#��֕���}^s���1GJ���p"㦊���/�5γ,�����,%����Xա+�'T�S������ "��ϛ7'����t)��<4�
����j�P���N���l�*`U�*�7�o���U�K ��_l�z�ͅʕ�uk�DJXt}����g��r�-]le����⩖?`$u���ѣFک��^�h���O��A�:�%@dt��_�!�Y2��z�菶�sV��o����r��҃H���߾p��6�l��K���ucM��7�;�X{�7m�;o��X�1�j���9~cepek鏚<�C{����I'��qEz��ɖ�����X<idۺ�
�q����D��5���6��E�16+N��)�ڳW?w|Ѩ,��ұ8۝�G�qd�%h��/nuI���������1�!X�����`@�����EX3��T�9�����v����g��΀uk�\x��fw�����������l���L�GڅDR�IEwmIG��3jC� ���`+�k�[k4��ZUB_h�x�-F��z���3�XU7ը�t4(��q���ϱa1G��F����u5��M�t������0�Q��ţ�������hL^עB;��3���|����ݖ�.�L��4`��UD}� k3�s�6�X�5�<�읩��\Եp3`͂���į~r5Vw�H �铞�e� �W��U/�BJ�r�6A����,,��*�zL1�~/�����n6ꘓ�!��(���֚r&<`�@j�#	����T؄�Ck#C��^��B;`��� ā$����R4ǅ#�o����#�����2�u��֢S6���B��M���葄����Lah����%Vee0��馔��hG�w��ń![��`���@y�y)k�b��6l��Lk�X�Ȉe֊wi�E���ģ���̭��6�3�=Z��֮��&�X��_X%^���p/�i]�]����]�l��+��dF�\����ՍaBˋ�V�Oe�z���C�\��#�V>��b�ʦ�Y�F<Kf
�m�Y�G(��5a0���W�WVg�8����͚�:ߟ�37��=l� ���7�{�f��QG+LJ�1V���ǍՕV�Kr ;W�~��w�]}�v��/�+oOF�°s����Y[ ����λ16�˿f� ɛ�kE�q{[&�b���2�XE+c�T�5��Je��L2X�X'-��S������ؒN�;hQΝ��,`j˛o�JR��K��t&i�p+c�F���I�@�f��d"2gN"�����<.L*�-�[u�0i!�^�z��ZV4�/��Y\�:��������y�d��5�ӧ���(`M�B�S�&�n�'�BO�����n����ZI:���{d���ԣEo�1��Pr��uG'��G��������
��t>Sm&���G1c�<����;�mݼ�����a�	����k�[�������η�uߨ������9��q�݆����^*xwV�g��D������DY�ݐ!��Gk] *	�ao��a�>*N<�|���^K�@�W?־��k<7�.��$�U!� �i{�td�F2�W��*̍�q}�k������oAR�B�Ů�Toæv����e�j��������ڵ�=\ �д �cMc�ۄ�!���^b��d?���[E-�/c�\�Yzm<�d����-����o3*8Xwdй�T� e��x�jT���'d���:o
SZ�+_����d%@� `R�4��7D�ȃ� �����^��+V�xi,�m2z���2VS�(48-Y��$�hi9]����
�zk�����g`X�n����\��Zx~�����LA��� ��߀iJ�d|�����'�s�*q}�z��sR����6T�lP���Ѽd�GɶE�x�U$h�W��/�ko0�D��n��S���-��}�,��B�R�+x�������L��R'h�M�H�}ZmX/ZS:�
~�v$b��dg\�r�{� BT�"�������u�{�K�>��'����R�.��6^��[�e���G *0MF��t �/��_���Ε �Ы�A�.y=İ�O%�`��9���M�(��2�:TJ�'�Q�/l��W�ZJs���1"O���"^��`�x��w����
���yɽlc-����2^�uue9-�M�5��:b?�򞷷ޝl���IC�X��'P�*H���~-U��g0����A���k"��^Wk}�#Ɵ��Q�R��j��n#�R*���_H#}�@��jc�Qg���&�h�K�UR�V!>�Kw;��,�A��P#g��VY1 j�&�X-5�V�F5�@�PY��$(�T��5Y�Mq�s�{�m`$�c�iŦr��r�h�i�8� ePiZ�$�>�z8���2P4N٭��t��\91�a������H5�#Y�>G�Xճ�PW�[�dR,������nZf�	Z�y9v��א����;K��w�,��B!���ݴ4����9d�m-�/>�uˍ$�K������c���L�Oz�^�4�-9%p��il\���j^���=��=	F��{mYG�^�R�;�M��7j	�=JL��*���	�Z�?f�X��=l��֫���t͵�4�`U���A��>��^S��������-]��V�k������L��0jѾy^>SY)�7���������X���&��U�|3c�R`�R��+K�C���N����y�ϳ�<��hȤ��!�u��� ۳O?��b{����7߰®Ŵ8B*�!i�T}�UzDL{��*8��e��Aoj�ݕ�g��D'a�i���)�ěB�F���V�#�&C��A�IX���i��o%Y�����DA�rD��Q�U�(eO��R�T�������?ɿӘKd��n�6�b�\J�$n�t�ۖ�%��t�V��;UJ}�,�>O��PmDdM<_��2�j�9Ұ*� 0������n�N����+����vP������+I��u�\j k�u��ENkz���5.N�\�T�K��OܰBm\�V�'���
WA�(ظ����ܶ�����4[�gϞΒ�c�<�]���=c��ũ�ZraO�X��X?�����7X�nU0������k���7p�����/�¦�nO�m!~���,r��� ->#�Q�$f?h�_�F�/C�`�����l0�C�����E���������5��%JW�!�j�|t�1�����_d󗭵�ߛm�i�0\Yٌ/C��V�;��=l�s�ňH�?t rq�N�M����t�]��tN���k�k#~�-$%-$Zue���/i�}�����m�)P��ۈ�]	����/O��ʞ�8�fL��
�:��̼"�Γ���V-�\�2V/�&�ʖٌ�t`ݚ*�1��Z��7����`��<�+�'I�T�uՈu�	v1�Qg��EԾ��F����*��v�&5��%����F��N���ӈЌ����і��z��Y��@����� H	��W�\J��e��cc��{?�V"�])�A7'��#�D�FC�.[��,FË$�I��(�KO�6�����I���҅���Ũe�,[m,\t�~��$�U�Y�2�-�QCr<�-ڱQC�9'��lQ?��[EY�ϴ�5�%JB��f��������v�{'���۔t+l�n#�%e�VM��Q�]�D�0�/AZtav�����	�kP'G�f�7��1�����zJw�'ok�u�2R�%%��'��O��7�y�O<�5�:h��^���K{3�=�{�}66�3w�gl��u>Y*�ָ�G����=w��-����-���L2�d�*��C;՚��<e�'no�%+��^5+;���I���f��_J��g�J���t�x���h�.�qGl��a���3Z.	��=���|J�U(�҈Z��W�v~�#hVfS�Z��+����6���}=/�z@$-�����Թ�^䉭���ލhf�!��E�[�}ϑQ����z÷�>�[�|���D��J����\DCգ��3�ce���`8}����[���ьkQ��_i�B�mm��	����g������y\�Bj��*��駜`�6Ʀ���^��:���%��˙]�`�O�},!��9�3����\�醵K��֊5�̊��o|����k+i���o�#�ŢG�bs����J6�rf� �s:��Y��6ZN,ǟMhO��h�d�p���=%M����;ei�}`���-77G��>�F�B���I�4�%jL#��k�,^��J7R���k�%��*
��!`$�A�?ƉS�$+�f Zjt�:sc�} �3`Y<��sR]D���
�ߪ����w)���V�i�J9\�&$+�/H}u���Hj��R�!}�bA6�����~}" ���wԣ��$��x�\��tc) ��d��"�Ǻ��8�UW]�c��n#~��S��52
��������Ll{�uJ� �	J��00
�J���O��\�>�,Z6�@]�ߠ�K'RҺ^���kV}���%����*x/�v�(>�_k�k$����qO��o���*�����1=�ze6g�2�p�B[�l��Z_f�N��NYH&i Vm~j���M^�+ V�Fs�U�Ԟ��c�F�0���S dKM�d�)� ;��ìW���:��&�k��R����ɝn���5��h���K
��T�2�}t׺�]b^D>ak7����?�'^|��Xk��]B���5��c� }����5|� �$M���6�*��\��D~ ����ʬ��&��5
Xr�;��c��#GY�յ �6T4{����'��/�bݻ�%�c���$���Ko���ǽ>e�=��D�.���6C���(��/@o\��6W�J�&e����O�~�LׯK�!�	�qfu�Q�Z���F[�d���w&Z���t�����!lմ�����[���L��NAk���+���u)Goni�}`���/�ki��+Ժ�����DE�7C���6�d�����7�8d��U0�՘�x�j|	�H%xiD0-d�T<	Q�J��
o�4�EI��)��4@3H���e�Gc16ъ6����x71GM�Z]�@����:�i���$�)=��J�gih��W3ǦE�I���{��{    IDAThc�j��uu�|��m����2��s����z	�d��m{����_n]���W�2VM�Qƚ���-݉�a�w�Zp�
e��]�cV��um��0�>P�![M�D��u�����U�h�"�ؙ�<��[�%e�'�t���-3V��$�"�N�ٙ��i?7V��K����Ֆ�jKm��^w�;WKۣ@hu�Y9��9L�,]n�UP�C�,akX�i�t's���jH�Z�X=��=��HJVֺ�l6t}f5��>�.:�4���0D�+|l�N�L���D��"�KL;i���'0��?U��,qS4�܍�� Z�����`�j��?�����k��8�K�Ld�n�&)MK�FI�� k��|��j�L5�ӡ���_ܒ��j�A�\ˤ0 R@�����
�d�ZB��\C-��ҡ�qα2��l����;}���� Hi�n���T�k�e��5����d���O��P��*c�<���>Cku�t͵WYo���k6�~�{T`��
t<�`__����Y��X?$QC\E�γ���b`��>�A��k�	����5I����u�W�c�q~Y*kU:�YK�/�R�D�`-�^�zY�>���K-X��'~T�i��c�ΙLD�ű���
RoT�覊R[�z%�k��bM5��4��;h =��y^=tBs9�jtL)��� I�:������Z"�6F)�\�f�-X��֮*�3��!C�#���|l�e0'o�%K�Y��nP}8�5Q�-@,��ĆI~3ϟ��[H�n:ѵ�$��8�æ�3��5)�
�Y�U�&�v�>���z�v�KT'f������c�OYY�n&������kS�]`;�>WQz߾}}й֐�J��%���X?m������e�h`{�Z' �=��������>��1��Tl��*PH�xe��^���s������J�zt�Ƞ ������&��TԝA�}Y�����s:��l�ɞ]��zؘ���� Qk��h�������9  ��0$@�CܔM��D�F=�����I ���U�XZ��շ�}�<Nv^a]{��}Qufup �{6���ͩ��XUނ*��v�	J5�Еj;lf�S0�D����U��!�6 ��]E ���ŵ)M�tB`d�6��z����i�Y�)(r͋X?V�������5�[��fXk6�|t����K3�٣�7��H}��6�U`�s�l�|�F�}�sf�g���ǝ획�kT�"��
�%`���-5�5L�	b��q�EHhx�jl\��%y-^��J4�����O���#�{���C�u��߮%;4�����4y{���a��<�2��������7�1� oK��9�������y�}��U�����3&�`���6k�\.^^���S}�}��A�>}�M���˿
��+�EU�g'T�����_{�������uԝ�m���٢�x^���F.қ�`�O��uV7v�LA��TlX/��J�XE��n���;j���������mS5�)��&f�!��EF����[�2�V	X����0�<vv�����w��XUc�1��y�Q�X��X�����#��*zT����T�0{iU[mo���ۏ�w��g�eM�X��߷سD������r�����m�=b��P�2P�fImx���E����ꡬ+_c}���5WЏ?�7b�f����J	,5M��ZP�"2O��+7ؔ�؂U��y����a-&+j�0/�zu�����A�ҽ 2��*+n&��k~� F�ZŞ0m�z��I�>{N�$ >�ڜP�A"N��D�%�XwX��E�f4T@'5��"U}D�vԒ���\oK�,)�_��z��6�E-BG/Z9UO�-��jU�?�%2�A���3��J����%�, �^������Wk%�:󥇬o�ȉ��&�:��!�?zl�ƚ�}��������oe�Î?�R�z��R;������$��
NK�`A�ʫ3�҅�o�F���+W��8e�z`��U�մᶫ���z����w��eD��s��d�}�Xɶ8�E9)��}�V,^��^���j#B9��=�X��]�������;x�]�����x�^~�+���H�s3)��a�"��n��V/[i�����
//����kq!���-Y���0~���Fb���s�3��s/X>\���põ���.@�W�5TٰA��;�]�d�}<�$���-C��OE���Ee4�D����븭�U��뮊�-�H��Jp�부3(r�5�%���V�$JXF��*�߲]'q=�ȿ�� ������"��#�?�W��#'�_�9�A���6�,��rjTe#�O�	q�bLi�����6t`�M~{��u����l��v���vЁx[���2��G?��M[���հ�K@��#�7M-x-�vS�&ֻо�������l� T#�^,�GpH}OY��{]y��5y�����u��wL�t�бI�H5\}�hR�Rǲ\��!b�w��9`8�(�2��l�T��R?�t^]t����-����1���6��Z�)!�� �2�OX���B'��k&���@����s`�րUl^>l�X	�֚jճS-�N�>��P�R�Q}��i���l��Ç�G��`����:}��D:�K���Bտ@�X�#�%,c�x�J_.��ؿ�J���x�%;�����tˍ'�<�ns��z�w~����4�����;�3V���/�q!;
�F�;l��[��~C;�j�X5�&
�`k�QVE����f���+l��e�����(���`}���O��Z���7l��o:�s��c��O����q�)�y����e�:mES������o��-[��n��6/X�¡����G�K~�5��ۨ1C�W�m���o�|�b��h%���=�{Zs�ԃ=�������{v�Zv!���-O��]Z�����^{���I ����������R��k��P��g�kH��hs@��-��$�<\�@���P[U�V�pqq1�;�WD���{z�q���3*X}�XE��Xw�L6��f��?�¼&�{�u$��R�XS�8�_7�0����_�?�q�u��ۆ���E0���G�g?�����GK�9� �c�����m�"̕U`�ܠ�%v��N����X!ɔ�Te~�ōȐ�Y����0�����+oؒ��ot�c�\p<2l�����Q��g�h��e�C'ˡ��چh�ؿ&3ƺQ~dx�SŭhC2�� �H��sW��/��/��t�E� �UV{{���O�
�#���Gm,u��E�P�I����J��A��.�)�A�J���=�v��H7�g��Ҁ`Mf/Y0i�=�*�����Gl��'o粞���v�+�'���xJeQ�Jd���U����#�48*�d�C�}Ձ���Zi{|�	gǾQ�{X�?�\;��lѢEv����j�[n��+Q��C؄5��Vن��Xs��O��^��KCQB%y����\f֬�{|��2�P�s���f�mw�o+5
�:rD?����m-�rV���"�.7l竴���x�I[�b�����3N=��+�m-���/�K�t	7B�{D�z��;�=�b���� 6���'m��X�9�4r�d�Wؤ�߳��8�y�L��V"9]� rIg��A'������sϷ�]����4�"di�>V�I�A�H�Q��+[�p-�Ps³���2�L���UFz��:e���f�	"�=�e+cU]��N��W���������ԙ�t�G�П��S��Z\+7C|�ab�D�u`�l���]e#�)��
[�z�u��ߺt��Cv�kt�o�����n[�������-�䀍������<���_�S違h�sP�O�o�td\Tsl������=ZER`�4�ʇ�;���1�t���2�A���$���瓽G�l<IL
;t� ��>�QCzZ�@��,���-/s�o?{�J�宇l��l��j��F�IǱ�Tp4ӹxb�qp�h�	�jGOm�2�L���)���m�'z)�v��� �lf.�N�.�p驾����S> ��f�� ���F�SQ��j��	(T2����u�m�K����.-.)�S
:�p���
�m�X 8����X�z(�M�5�w֨#O<߁U�WQ�{XE��5�c��6�B����`��>��g���M�i�J/���ˈ
�ӧ��[2o��WJ���Aė,��V�F;ڹ�.���R��B���,���l��e��;�*B��t�\
�Ǐf߼��������.�n$��gq˼��%�\��˰�[b��i������?8�t1�<y�=���d߫l��v���SK�k}��GQݣl5Ŧ/_IOl��d�Y��6�oO��߲�^}�z�)K��f�Di���*���B���j��^:����W��XKOw������XA�X%��S�2�4�(���K��]uU���S���!���54��5��f�V��*{�rW�d�y���{{C"�2n�h$��$�֤L�y�����	�^U���O��Z�-�GT�zI�����~�m�}z�!#ڡ��A�E��}Ѥ��j���뙹��f�]`+וۆ�j�)6`����3�,UkFb�T�v)A�y0� 7zhDĒ��E����Z]_��n��#(Vs�P�"#7�,���irk�X�%imf"�l��'�2x]�k��L�5+jД	�Vm$[N��/=��6�(�B��E��j�@i�~#A�OM��y�Z����wAMȮ"5����XU� ��\�=	�b�E�f�PK�����H�ę@�*ݛ
������0��(@H˄U`X�wSp-j�Nn��)^�k�\*��ԅ�ڻ@��\��P�(� ����t`-)���z��E����C�u[�%G���w1�،Y���TǠs���Vc�#���~�����2���
�tѪʄ�f�hL�X+4�A�����&�.^�� ֱ�I�t�m�@V?�7��-۰�b�ߟf�k;�ر֯w����=7�:���i���?t��ڳ���s�S��D}~òɧb��޵��'-UP:DS��UVVA�S�)��=���#Ȍ߳G��u�A��o����I{��W۩`�X!m��j:�b�6�ZK�FK��;�]<��{�Q���S��Z���F�aʽ�FEl���j�M�c��
�ZA==��ܬݻw'J���\R���ɠ�@�+�	�<@~}b��D�>\��&�l{t��/�su��
{���3}n(�Tn�
,�3�(X���u/���	���U^��*����M١�n��vܘB�ԖRWۺ����<�Y���.Ye3E�j�܋�T�$ӸǤ��'�Ө �l~^�����u����f@��k�F
5K�u=�V=/���v��Z%������$3��G�Eճde9dZ��Ҫ}��E��j9���h&st�V�L��L-9�!#W�;�N��(�W��eJ�^EX�D��J�����g.��"JLW>�.�
F3�\cP�qj���!+Q&��� ]����kY:^e�$>rVjlS �=��ڲ����!��l�W � E�'�Y�7�ZϢ\+��_M;G}� ٰs��q�1p`��
`��,&�P��z��y�Y0 b����R��o���:�J$22i�b�j ����LW���Q'_��u�6[V9/�����<e�����OY��T�kN��S�*X궅�x鐓�B�:�6�Q��է[���o�¹��W���`{���i�Rد���o�۫����9N:� ���S�T�/a�_PT�c.���4�������m�����x�/� T����c�����R��>}��s��P����M��_|	q��0��jU+�f��GK�T=�C��g������?���3zZ7q�_�DNn`!5 ��� Ve�X5�&d��sk+c�(� ц_PO�m'c��5��
XN��`�^jo����jg5��:��NY���t��D��]ݟM�(8d�ʶ���w:�r�J"�� ���
.o�T�{��w������ݓ�hј��M�.�beY���������][���Kl.A�J�U�l�6N�Z2١Zv�N4�M�9b����ݭ��>�z�W^d�9�`�M��X�K͓�>��<��އm9}4�ݨ��VUjV��$o��3���U*be�Q;�� ��)�t��7OuQ֪���G�ך7a˗�d7\v��|�0C��@ő�6JH�V?~6������<���=2@ў�CGk���i���L&� �1d����87����{�{*�Z'����٣�?�0;p�����l6�,Rj�r��1��fw/ʱ3O>�[o��!w\ʢ6.�u!�����^ۊJK9��չښ�t^S�̤��!<�1s�=��ì�ʏ���9�� B{����}zZ�����m�ݤ'P�[��w.c�
�J��%�y��1��y����]w���n��m���s������Yْ��=cM��=p�i���Dh$�;��|�*[�����މ�Dn�+$�������������'�w�+O�ū�l�T�rT��K~�_iO��Q����ПD�9g�l@f�l ��Qc��ߥv�]��}�ژ1�\�ha���r,+W^�x�b�E��^x�-+�	&��W�[;��u��b�G�`H����.�MD����9�X��j?HW�P�R�h#��l�����Z1j,o�>J\�-Զl����l���A���O�6=z��(3�_w���|��+���wt��l&�hl[)����m�Xkˣ�������%�0�Ƃ������0�$�Α�}��3T��� �Q��4����8��#mk�f��,����j4JTd�^���L6|��4 �����FI�z[T���N�e#=�ǌb?�֥��P�˝��XM���sV���~�g�p�Z+�?�2署�v"�1�
X��DY�� �6=���J6Z.k�"��G��9�l�69C楶X�#�RO��W�~=��u� '�'+�z�̵��ͷ?boM�g��l�����K�6b�¨�8�N�"��+� ��{��J_��*ߋc��Y��P�`���Gn��i�sm��o��f�[b�9��4��^���	�~������es�W�M��m�+'32�@	��l!X՗�By0Y5s���J��/	X�4���!
l͚�z��:YBF߫]T��H%$N��CY7D�U�PΚ7�l%�N���X�	�1,�`��9s�G�h;�$���&dNj�(-]絸�X�m�K�`q�O����Q���S��'����bp�s��	ݓ����.��g��YC�=��֋v�cyn���j�?c�u����Ioa�Ua�bC���v78� BSc�._����|*�'Y�>���C�l"�(��Q�[�M��K��W��״��u�LY(��;�3ޙ��˹Cǡ�蚠�@D��)�hL����`�X%aOC�(U�g�P�RR���B;��\���?��({	�<h��� �I��Q[�8��kC�)��G�6�zW6��@3�sB��Z#���Uk~��=cU�U��6����;W��{��f��Z֐�d@�J��%�@��y��%�g���H'K�yM3٣�"'��}a5�s�r��B0�5~jx�4 .����ǌd~h��:��eX91ح�?g�<���� rX��7މ���m��^�6����48@`$us2z�#�a ��V��U�K���v5�C]��k��㏲k.:͊%<�=�ӽ���m��'͵��~?&t.�+Д�]��\����>��6%>������29Ɓ��W���!N�uv��rR���)�I>�͸C��ǎ�_��^[�z�a�B�����Kh���K���:
n��7�Ƹ�Y����b4��&�ځU�K)���X?x`�^�5V:Ч�!s��S�ZP'R��C��L����u�+%�J0b�|:�
X��5K�-�U&���.8�9�=�L�Lt�	?��	����%Ly@���k�E���J:��%�^h�t��'�U�)�P������In$J�{J�7a��?�j��x+
�t}�G�B���+97k&
V��ld��P�6�j[[�|a�%�Z+��ߚ�H�\�2<up    IDAT���9���i0�JӤ����L�&�Cs�yLoM��l۝Vx�j�t.*X�*���T���)��jӑ�B�ZM�@4��F�)����� T�6��}н��(�]ݞ#r�$�K�C-BV�G}�f�jx�nDm��56����w뮞�O�uVQ��I�TO��?ea�G��������V0�8>Jf(n	P3A�4�	�^�)+��^}k���%et�_��ʭoa������޴e�(&r`j��j�~~oA���o�l��H�i�Aې�		����A@��D��P�Fm��^L@\�w-ْ�\[Da�\�S�����5V��l��&�RB�A	�b��uQ��~�>�^�.�$�ƛ~�BX�����g׀U�4 ��!�qw���Q�_]�Cȃƌ����wߵ���p~7U��9q���M|�����S��j\�<������7�{�ޟ1�Z���PdkJ������^�o��������wVZ�,ʘ��5��L�`�'+c��B%X�}�+�KL�ܧG//�Pڙm��n��j޺եkW��z:C!*c�/��^��-^����1Q�y��n�}��/��*Pe����j{�F�5`��R��p�B{�W��ۈ*��O�i��h��#�x^*����j�\Dd���Ϫ� �"	�
�`��0�F�H�ӥ�k�\]tOd��m��@���VM͐��j٩��Pە䝾�L��d���M���]���J ^���,�SYhUPg��/��٬
 ɸ"�6ܜ�&���'O�GFۮ��a�Avf��j�V��h�)xH!��#�<$^� ��f���m	�qَn�>���t�<x�-�D�Mp��q�UHA��'��LѨ@]��>V���'(�'�ތuG���<��*�Ro�a���7l�]{�wH���l^�؈�hO�U���@��#�?>h�g�vĪzW6�uV�񇌰�q�u��y�ER����@�n�5��ɗ-��j��ئ6jD�}.���8%���/��2O6�)'g_����YҌ�������LX��D]��٠�)2��>"ʸ�F=�WKm��v�!���N�BRJ�Y��U$�0U���>{e�l-h�wX�CA5���z<�v�� մ&s�av��'ٛ�&;�:v�~��So�3O?�L�eW^a�����"�R�7�r�:;�qv�9G�o���A�`5�s�����֨^��~��o�{���_[%�\�����i�&؈`��X��N}�Q��R+$��ꛗ[ߞ�X��n��J�=E������>�����K�:��C�k*��G�� �����3�e��6��\F���{�ƥ���R�)�J��~h`}�-7{eU�ds����Ǡ��C�}B঒uQ��fU*���G��nZ��,\��"���T~�ٌ��
Ǥ��/���*��*r�t��4�[�M7�L��Bt7XCm$�Ne�k-�t
2xE]ʎ=�ujHv^Q[�z��u��+	>Ѩ�L����-V��n�Ųi��8�༔�qq{��j�&�N�Q┐D;-þ�ʲs��eGL��h��Z�b�6�;����Z~1��cg �`ѿ�X���C��{Є_kL�=r�H��GB��� \�fم>�\f]j�L����ڷ��8���d1�����9�VG��2+�G��	 �k#�lE�?	F��ɫAJ��5����������+:j�R�6�-�Ng�<��A�W/���ւ]?��}��G�-�KO�����>�EI�t'�iWƲ� v��\[��.��,;���������؟�����3+w�f���aۂ3����21��TC/(��hd�$���~����b��M�7��v�#��{�ZzC�*C��hiX�1�o���T����mX#&At)���^��˼���_��l���_�@t6=�ո�q� ��C/�k��t2�@�}��'O8�0�⢣�׿~�&O�n�Ž��Dы�I�?�ݵ�톫� Hγ_p�(õ��J ������ٴR�r�U��%�o*#c�x?IG���t���?o��}4� d�:��^�c��~
�f8�J��H��.\���>�=���t��L�iXe�MϒV�}��c�DU7�է�f����@�rl�u��Y�&�@	��6j�����D�&�]�~����r5���X�I�p9�.��UCRo.�L��ޡ�Q6��xTh�@<��N�.�E#v	û[�h��h*}���2��D�r��谉�Mnj\DK������� A}l|���Kf/E"t�p;)����ƂHa���w������^('E���Q�Hc�G�S,��v���q�%Q��}��I~�4�F7ӎ���ֶ* �uS&(7�0@!L���V1غz1���3]C�����N�ݝ-=4��=t��M�0�?[k��_�<������n��5�bo���O�tb��0�f
�ç�d�i����8����ۇ�qMc��̓\��.<�DD�Ŷn}�����֘�J�u��~v�	{O����'��
���.LGA�P�ծ�.?�Lp�[j{u�%1?l֓��Oo�ϖ��ԥ;�3{ϓ(��������m�½�R�֮>�D�p�ب'��᱗��o���x������N@�ʼ�݀��]��M�"�W�zmE�&�������C֦�V�Ƀj�R<5i�����&��{z?�eF��"��8W߹��>�G��̠so���=Ծ�=��S�~\	t�j�Gy�+�gL��um�B_:�$�4/��i��2s��P�dO�._o����]}�i�ӟ�eSg��s+�t��	Xjʬ���#������?�����Y�iY�����a�a��T�PT�;QQ��\�u���o������؅��*b �Hw3�t��{�����Y)׏/�~\`�;~�w��\���������z�Ce�̕�?k?�"T�
�>UpE@_~��ֹc'Fmf{�ZJ���؏�7+��
*o����9�� �K>O%���`DH�!�%�i��yl����%7����7m��P��_��� �Z�?�>@Xg�?��|�a�������X<�����)�5�J���	�8�ݚ�R�
R�YF����ٹ/�ke�ޡ�[ң�ޝ~7�ݎv2!Ŭ�]ﷂ�!U2a�S�h����TU���鹆R��} �I��T�����y7}��U7���Nt�*V��Ҹ++�+�q�QTc�q5J �@���ۆ@A����X�tk�����kK��c�g'�^z��n¯9V屾�����&R�nA���%2��9�1�W}�ДA�n�t�u�C0U����e��;[z���hi����6�~6�	Xt��8�F*�]s��s�w��ja��Gs�q�l�UUp��y�<�E���EU5a�=ڶ���|����ٝ�~��;�6��:�߉$��|�H�������x��G
 �I�η[.?ˎ���O��H���:h��笱��=�6�RA!��'ծ_����rd1���8�PEv�������r'(�>��G��'^��E8�*���^O�`��A��'�.*W�9��Xf���";d�6�D���c}��|yk�"�������o���ym��� ֛����Xt��Yk����qF`g��[�Qj"��MF3b������x�o���*�omt=�ϘC�&�cw���m�����U���XQ�Xi���$Τmw��g�)��#O�>���|��I��Isw{Zk��l��3_k�l�Z2�x���Y��]lk(^
��ق�+[���b:`�>�**X��mb ԁǝ�s��}`��U������`�;܁l޼y�A)��7��UL�� �GϽ|�"�C4H��٠a�Y �c��T�	8�)x�]���Ţ^tnP%����՞n��`H�Z2Q=J��Mpscg��A�Lp��I�h�?R���h��N:��S�
1��
�NsA	�w6����U^�!��&�ފ5��fX����J_���>���m�JD�p�*3l�%Z�/`Ո��m�zx���e�Xw���#��#dzT�8��޹���J�TY
">�cP���v������ ����k��_���c����n�87"����!��x�%��k�s8���U�ٰ��������)]T{k�r��ݏZ5b�*ZP����a��*�gW�Ry
X�� #��f�Qv�у�Q�9浏���&XMz[6�2K�� �6�Gy�0�w<�!��n�-�ߨ�֡=���Z�U�ϳ~0}����ɬ���)`U1�
f=���X���,�����x~C��ә�DX$9�%Ȉ�����x�=���ni�S�����ߵ�~A0I,`�]�gl�R��C,X�-_U���ӞǪ<�Z� %��XŢB�O���^6c�zź`�<VgP#>��ݦ�|�,��G�һ7Ѡ��43�9�J.��v�=�f�V���P��4��R�\����S.r�ޟ���Ox�B�h8��������X��hk��l�m{2����K�KE��F�����=(IA
ݰ���O�䒢�G4�v@�'$��7�~�z'�KU8��5��Z�>2��*�������E�юD�Z��<� |'V��F]�����X��O�ȁU�q��[/miY�QtE�hx�����4�k4�#�5�o�%:��Rռ�<ְb��[:����&�@%�k�_O�MS0u���nӪ��8�82��a�����ˤ�m�GSh�d���e�`^�-���=@`x=V����*p,[k���B;j�Ό���l�L�ۼ|o�Z��ݏXmj`Y�"R��� !̙7�f�=��U��k�9�F7�����?�{ǎ���qNb�H��*W����@�G��K*<],W�ֶ��+ε����U�����dm$mg�+�O�<je񙬁L,DktŪ��wU�[V�kZkj�iz���00?e[KǢ�F�T��X�r[fZ6�y
9��dpR,�m1�B)�:�t$�Њc#�)O���0�)��DK��#3M���E�o�W�b�`�T��\;��<_�x�M�8�ۂ�b_��#�&`6�k�#�q ��Td-�K����������9��Pt�5	>y֤׬,��uv�W��/�L�p�&e���%���4;�he�k�f�P@*?���X���d��y�m+G̔��� �K�4��)P�̻�l;��İ�KIe�)J~�^M~ɲ5�#�!��	 Q:��
V���$���X���7�2~�n6�Q%�+�E��(a���}(�EY�9�i��ݵn��E_~��&`�sX�����M[�4����|$&�hC���A4����i�[z����:�+V��v�O���6�������]��5G�����Ҷ����@&�{/�{�e��C���#N�ι2�S���¯W��vL�V.�Ch�yf�OlƢu����زb@E�FpD7�o\K��LqH/l�7�ְ�Ŧ����U���c�4�
Xi�G�\��r�,\m�F�����T�ٳo}e��y���5·:�*�wͶz�̴�z����B�e�U�o���wJ��9��F�/����۝��ڴ|�'���S�4T����X7]��3�z�ڨ����n��4j��a��V��n��b9UN�_wMc.���Zv����Ĩ�백�VC��<r����Jb�X���yH��˩`h�|���<V�$���*k�51�)�zh�Ut�c�͘�M�9í$wz�[kXW�**X�%���<����}�����w`Ѫ��^����T��-�q:h�̷5��޳;٠�O��6=�eJ.���0ۓC�x��j��[?�}�e0��c�O�.p!G|=��{/;�ࡸ#qAS�
�˰�z�Og�ǯ�5�p*�9�����Ȍ<h%L�*!�/#��8�z���ɟ1�J�,|. ͔�l`���U��RV�uGQ��ADs��0���h��a�B4�F���W}-E���:���t�X� ������/;V�2m �R�S���q�����=�}��'،������8�t�����Q7	̖�������{�,kH��3�m�VW���#�ӆ�0�ժGuL�K��
��w�}<k�e���z�6�n<��'BG�AkR�'���r;���8�L䨍{k�=���u����C���4�ӨD6� ��7��"UE�_�<��mWZ[�P g�� ��{�s��W&Z.c�cm���|�U;Xu��c�O	&A����/T�(?b�/� BJ���E�!��6�c]�|G ,�3P	5w�-���g���`��+j���?�y���yv�g[N6T>�Sz/�h~�j���n�h����	oX!�8��9���S�J����g�c{ｷ[
X5_��٘E�!�������%���\���E�w�I������l��e�����~�]��:��m��"{��bf�d�Ņ��Ȍ� ��?��|�<�b��,��9�v�IGe�����cm1q��m���W���ʐ�)M!FrY%�o/���#m��۸��w�ae���nDԼ�*�+����KR+�U�%�R����J5`�jh.��ԯ��#��hn�;ۺ��ϯ��S'ԟ��O�]�GS>h�]=�m=����k`|N�N���VU����u�������ͷg��*~^,JYhS	P=���m���}tF�կ���l6&�ÓZ0���"u<�VU\`���|�%�Y'� t��YKo^�S%���>�Ǟ{�� �8z��0�q=��PU�?�Ҍ ���hSu�ʹN�[ Gŵ"���ֵ x@Es�>8�֚����9��
Unq��ҳ=�����Y��(dD�Z�����l��~��*�It�[���u�{��5!�>��U���%y&+H$���G��AiԴ�V4���-�-�K-���_�D_	l����H����*�����h*D�*yQ���T�^��XW��	OZc	Ǚ��L��W~_�"���F��vVNbS>�z��`Ht��a��n�����U�j*�CU��*V,X��~�a�
A5lr�TB�Y�N��m:P-j�!����ew��걶�������`����K����]���h�#&�7���-q#��(�V} s2��)-.b�WܚV.���;�����^'��;�����Q�ؽ���}����xz	��PL��n�����d2�F5���N�K.���X�U�V	�D�li�uKKf�PXy6���7K�@�+��:d)B�ݒ%��_�t��$^�J���hn�xiKG���}����I�����%1��-|��gp��%�|"Y��ަ��G-76���=Ԩ�Àa����Ϡ�T��#0`V������˵ۮ�����a�G�C)����n�?�/�K�zp^�F��/�#;ZI��4Y���
��+��g"&1��SR�-���e�P�Y4���CcE�2���Fِ��3~�W�,����^R`���kK�1R�����v����vBi�{Ф�[�� ��0E#��l����@$A��,�4U>é:ld�/	�Q�t��b���Q�i{1K�6¯�
f$*"^����و��F�A����5�ɿ�_  ڼ��/D����k}DU�FJb&�6%1]��#w@ź`U�UœKؼ	X�9VQ�g��)6���i���p���LbǶ�G����c��2�[_"R;�n�q��Z��i�k+��:�ϳ���[�.]��7&��O>�\ Z����z�&��P������S��ѹ����;�__��ګoO��6����7]�T���[6@�i���w�k�i�?�i9�--�M � Q�������{�ځ��i>ns�c�����Sz�Ӱy�(���[�Dz��_}���:�!s��t�4�ZÎ-Y��� �ǻ�~�w����t��s��OX���w�ͱ���j5�������d�	��?�?�O����q���$��({����J�#P9)�ʆPv��sM�$HP�2| h���s�a�J���{R���6�u�\`�鎳$��y�p��M|)k�}c_���(0���)��J%�R�2S��x�m��w�YD ��M�l�~F��q%��}��Wږ��5#�e������v�#�k���$���pl"c������O�L2�YM;�olN見U�b����̊�Fg    IDAT{>�����
Tt�2�>�
�'�qQ���<Uq.�0~��\l�jb~G�+k?+��D����
6�Z�6�/?������)���Rx@`ۼb���?"�&��h܋�M��t�7vo��]=�u�U����
^�l�	Xe�Gh���救~�nݼ�\���wC1�z�����PW�cM梯�.C)��
��#���V�H�e���/�i�V��
�ƣXKd�I��U�����Q͒��"�=�t#M� (�\W�>��������9�(��z؁vƙG���|ʦ�X���%�nmڷ����߮h�冕F/k�Y(J[��U�K��+�|��/,-Sr��'T���d¯cZ�\��bDyl�*��X@��5��~x��f�}��'ݬ�7�%�z���ɩK=�td���ЋR��J�ٞÿSׁ�RC h�/z5�p	 50:�l�ݻtx* "@��e��j # T@��m�P�v
X7����أ�IWL� G�&{ъ�|ۻ�nv����4.=���JO`�i�/`����_]l-�u��ba���e�.]�[*-b��=\MX�)y�0�U6�~F����m��f��s^����3�-��^�E�؋
٦�,՘M���M���+��~lYm;{���og���>󯑚�Q���*z��-��5�GC'�M�"NOuE��{�igM��?��y�u\����Ϋ�m�')�D�a7Kt�N�o�>��ј�ރW�[/��w�6�E��U������ k���I�qˑl8��DZ��M;��;'l��= �
�>��U=V��=V=y4�M�{Z �m��T1.`ց�eg��RB��V&��+9���_�223 �a���=��-��o̳/�*^bi���4�u����5�e-�������r�5�v���v�	�ؿo����&��~ǯl՚���_������~���m�[S�g_�,�*�C�3��:۵��m鱆�L% ���%ni��x#��^�_�K"��NZ6��n�����W�SW����L�����>Rr�aoD*�؄t�TZ��'�J!�%���pv�Sh1F���&eч�B�6GL��x_y��g_uO���d�#ĺ� �2��-�k��u�M[�tBf+j����fcs�nu�7��EU����t�#��P����؃ό����U�"Z�EkV���ygZA?�b��.��M�(�HR=�ب�8	]���@-W�
i^�V�����U�n���H��)0�"K	�s�����\k�ףTטI��hs����5\��k'��2��U�����n� J_�%���P�s����\z��Q4��=��V����+�����)`�`&8&�/��q�:u��g�f��7���oz}������q�xs�z�%Q�U_#����ֈ�v8�J��@V�u�Լ�M	렋
n�KX����%�z��@�l/�TB@�}*��$n�*.�LFkV,�o'�|�]}�p�������%#���FQR3ZJ�wCxѱ�Ӹ)֬\b{�k�������E��#c,k�j��O=�8zx�헷�O� ;��}����
�Q�%�'Z����6̮fw���-8/��h`�=�yI���;'Wy�)�X��e�	`&����/�E�%�&�����0�|K�6;mM��8��J��]�6q�~��5=�Zb�ʘ���:��2�W�8�좂�ӵ/%�J���hEy�∯#`�t��ڿ�+S07@�.��		`�S}R(����(������M[�ђ�1�Bgj�q��jU+2�gG��gZ7�c�T�	��|w C;�S>��4��Fx���cʧW�Rhf���D�S	pKݫ�����B��G���!%A��3�x�V�X�e}���S���&AK,m�*^I0�]}����>���i���r���a�O�t�XU�|^1!�J��4���Dī�I~F1��$JX�6�%EȽ�ǉt�w60���T�'<��m�Z�k��5n3�ub������0RϚ5�P���z��k�	z��*8�͍z���eiX;�À���<f���X�<c���(�MnE$���$ES��#7���(yyA(�R�z��(�"\�kJ�^V�$ݍ�[�K����+=Ѧ��2���/��x��ǿ�EK�y ���-�h�_��p*'s�}����Y!�!V~bF�:��޿�fm��3 \�O�[Z���/n�:�^@F�}>c6. OXN^Gz�A����5֣�GVe[���ll�4l�'$`Mn��~+�v��&��mE^��U�o5���Ol�V�r?��H*i��"Bɴ�� �j�A�Ɛ�Q��I/���/���Gyre��@��2K���DJ�TCv�U��A{��J���Ͻn����B���a����<\c:�~���l�����I�t�:�6Y�����㨦�DbȊ�쒑���'q:8A��0@b7Ti����|m��9����(�?��<aN��F%�(Hek��R� �-*xhsqC���d�xˀ�LѲ���hg�Gzʑ�|fU�8o�=y5�-�������g�[C
�Z<�E��g�s�5T���n��.ŊT�Ag|.-�Zz��q���0�y�����o��|���u��J]l�"?Ֆ<�?k[����ڔ���ya#��,e������u\4�D�?�ظ5�yY�nӫGO�&��{�������$^�d���ǚ̚޵[g�q-�����\�n#���c���5`����z�9�#���"$^
s?�@p �ʵ)�T�4�'��Vp�.XK�+�����Ұ����;�W_�:�kx�
��)�o��(�3O�l3g�r{�,����J*K���k����C�+/��,C�U�I�w�ܜ{m�g�2�j*�DT|�]+����N�����x��Gl��U�&��(+���\�8�(������|�us���U=ւ��؁C�҉�&�D\�2�Pй����t��\P��Mia�����zЬ��G��@7;�q�X��Г��du,>edbۊ��������"�7����}Ә���WB(��P��l-�K�������$ͥV*-�1*�xX���K�֋ϰ�N:��R�;�1�>�W��Ax���5��h���6+�.;s�5��Ɉ5V}=	/ *7��$_���U6��W�["5T�x�Q�f[���a��:-�ד�����.�b���)����T U�T6�k��z���w�>�ȩ���,1l$��|i��%v'��012�I"�C׽3U܎��TtJ�Q��#0%��	�_0�G�"�gE�@ˮ�O;Ĥ�Y��4���ϡ�z�>����Q���j��<ܙ���|ג|�A�ֹ���KP�{�ѱT�T�,�ut���B���B���]܁T�s�;�5;�-p��'vm��P{ny���ò`5n3k�Wt�:�_�P�!Pm�ɇ4^h�'>;[�;}5g��\�̾�r�)�B�KDdt�+��b@�m��Z��#Ρ�X�a��u���h�G�ȡ�Z3�*�b��U� n�s�v֮m��O���\�b5	V�@
��� o^v��i�����|��+$'�� 5�F}�(�s]���wk�c��4�,k���^�JM(�����vn�jOb�1��k;M��t+_0T$jW, -�) VT���K�TD�;�c��C��b�ʣ����3�n�;�� �t���b�٨�l�~ݭ�H�[��O����b2;�V&Z&z�
W��Pj��۷��,�����U��0�HD�������Xص0oܰ
��6
��}��jM���M�ěj�aiS���g^|����S<n3-b�����Mʝ
ֱ�M7�G�O�����L�d��l犒Bk���^�:��gsS|����+U�!TY7�[Yb�׃�|C	���`f�]d4��[2��`7����N��O{�%�x=��k����0��H ��Ɵ_@���y%b��ҋ��<���K�ϙnC�?��=�x{��)��o�rC�\kĹ/N"2Ο�hu~۸�".��7��*ݦ������m�6�R�'`��T�z�����ϭ��Ίu��wN̯��ok��c�>����|w�g8˨7�ex�@ �	�g�d��3gڧ�|�� F�Q��Nv�,L�`
���hH��,ю� ��Ż잋ګ� �&�^����X&ߔ��Kfw+��z$ �[l��CI�㒞��:>�3&��%׻_&>�쪥Z���R�-� YF�=VU�����yBN����c]�h�����JfI�H#%]�����oF��㰽&�?�R�u��s��
U@*չ6pa���U�ʄ_����9u#Up"=�zW.���p?�W�<��2��@3Y��u��Gbl����3��C����	��`�@eԈ�rņ�e��:ǲA�e�����T�f @�k!�$�C��
�QהX�����ΰ!��H�3��*�
*S�IA����_ƿ3͞�-[��
6��z�H� ��;�ʙ���
M�jM%�w�#zwik'uc5�]��~���jm���\�5�P�}��������RB�� �kŘ1ӪW�ek�`Q�n-�,6nSz\d>7�#m]	��MO+���LE���HqQE�Wk�D���e�#)|��e�O�Q��.8������\�L�����2��[�����C�O�E�Ԙ����~fӿ\e�>��+Ϫj�ɛܩ`
��6ss���~�����ۦO�fOо�H��W�2��/}�=�^屶��q`�|�tڂ���.M�q�6�i�Fr�E�n����w����9qmU ��#:}q�P�A
i6��%6{��VƬeԥ��k�����JC,\ ����[M%��d��U���Q�ZZ��ni(�D}�ɋ����7;#�j��f�����4���o�X���d���U�^�*��\t̜��th��H:�`�"�#(D�mj���T�+���A�TRɅ�q`��c]���̱���|OX�����mVf*`�Y=X>�6$��S�d��&M����.^�9��nU׵�?=���QA����R�sl}e�eu�V%gQU�ԗ��m~8���W
�m"�h��YHk`��*Jmp����η<���}��L���뺵�T�,�7�_w;��6�������S/[m"�U��k<�f�=��\%ה���a��
,M�ݭU�pH�M�D�$7ա�)�Vۓ/O�i�W�q<��6�����=jO����^�U�_g'��?�k��hi����5����9�U#�'F�Z�-\ow>�$�� {k`x�FT�*$�Ы~qC�%�
Vvmtl\�����U�P�����]�9йQ���O?����{�$��6v�X�d��1�6l������b"�Ԃ]�q��tȞv���~��,X����S���њ��l�l�O�l�yg��c���[�`��?ݡJ�w�h6 w&��uK�+8/)ݦ��s�xйz��>�\�:?¬�ҶQ[��Y.8Kl���1���4�B��*�\U�2.�9\�� �g��/��(`M"px�dL�#�f�6��6�V��ҍ%��)��e��l�rO��N��B�@е3$-���:��ڀ���R���Fm�$p���K�/���^�g=��#�a�Ĉ��V�	M?i���O`�Y�������7�x5��&`�SL��	#T��5��>�*�V9y�~+<�o��8V�~#=֟z�* � ��;w�}���gYu�{�{���]�T�H�T��Q�.$�*�m��w����Wk��%A�J�F��ܣq2��9��#��ZJ;A �%+�eKK&�r9�h�i�����ۢ����V�f5ʁCw���[7A��o����k�l;��c툡�a��q"�'��e��k`�Y�����߳w�ΰ��J,݃�����_�w�c��f��]}�Av։��]�]0���Uͬy^�5��$!a�*�������߶ep�u��5��
|5O�QZ3��W��=����S�=���o ���k`V��������g�����n������9�L���jI�]�uG� ���|:�0�A5X�x�nv�����z�f�[���g���le?��
�4O�'�sQh
kxa(7�t��a���C����8�*���R&��jz��_�k�[�\z�u�4H�*��(EQP��~��A�٣��Xt>g�<<H�i��{n��8H7��t����5XS�I�3&tV?�)yt~��)G�3Ѡ�ۛ�~���t
���?b�%w�����+^�'{E���K��B�.�*$��tqaj������jU)N1�[Qo��F@#�������Q���54���1˗�j"��6��1��Nj�t��"�E�'�cAUגF��w�a��˯fٓ�<���*P��T����h�.U��\�?��J� �Y�8�ܫj�h��С�u�w�|� <���c)g=��;M�r�=It���x�gS9U��oc��g�GS0"4�ڑHJ�&ʰCL#�������n���X�
T_�e*1��T�<O��3�)6s�*���\g�JJ�n����b�.�㏴�{tu�T>�ל��d�!�)�%5-�#G~n����2b�G��:V3�b��o�����n�����g��\�>��kh��׷��s��'�8+�cv��׸y�NT5B���|��.Zb�T����nQX�z��<v_;c�Q��;���DP��ۆ]ڦ����/��c��Zf�V�[��1���_�n�篢U���z�z?�j�,��L^�k��mbV�������|i�>J�^���m=V}[�����k9-�y�:��v�e}�s�U�9�k���-�X㨰T9��Zh|z{�|ĵ#�w
��CJX=Te	��5��G�⥴n�] ��Ů���@P�bn|�1�Oh��Z\u����/F.��Z���x"_�cg)���� �#)5ۺ��`�*8����A�W���
��z�7�ۈv�^��m��?��׍�#ݐ�Xe���T9�&�g/�B�HR�U���o���ڢ莗�L���]=��|m��5#m�CR�9�ʆ��є~"*��ʷ��t˵�dݺv�Z���M4�l6��9���/�Es��)*�*֒x*=6-��W$�ܿ��I�(��fe��h{��l�1�ӿk���y4U��#�<T���]�#�;S�لw?�PԊ�Ԇ�/b�c�����A�]���Vj]�y�>��M�&����R{��%�*��n����@Uň���z���������PI�neeKl-����R�	�qԽ��3�굫��p��k`9�q�{��z����o���>�1eunWXb������9����V�نr\�ۧ?ֲ���M�qo�c)Y-�����Uݢa�5����z�̱^|��ֳ{�={��X�I?���>}[�\X[�e *��ysQkܦ��g�&��wh��d���*�
l���ݷUܗ_~��mg���D���_��1�$cؚ�b�*[��6z��aZ�=�Tn^���|ye'�[�EVfΞhU��x���[f
��Й�Q#;�\U(%�� �2$4���{���V-�I'f�
��D�bM*X�`kNv�]y���)�%y���{��CM&-l(~ʏp�F�Z=�v��9�j�.���X�h�\��ѱ#��
��Fk��h/��)2�����`�����c|Jg]2�ge�K�?���^����G��&;�j�qTBQ��|	T^5�VK݊�8�!4�i�R`��`�>��ej���|��t���z��v��ݍ���"�J宬��+,�M�*��56��Y�|�:�ӧ��GwK�������	���B�&��N,���5E�6��I�ڻYa5/D��z��y�O��_�`}^�0h�VLb }R�d�H���aflSe�Ւu�ѧ��<��*��ė'��mBӟ�̊���[2���|ǈ�gǖ6tP+h�u�`�Z���x�R�(^o{�ݮ�lk�}0e�eq?u�DGUv�}��~��[��z}�[�c�Mu:Tpպ�6��'�&Zky����;v�i�>�^xO���X�C�f2m²b��/�b<[w�F�u�����"0��K��**8�X�������sY���~
�=�+א��<��;B�X�ѳ�"E�h0����    IDAT���A�b�ZP���0V�C;�R�\.	�j���͢�JQo��\U��!9(k%�����ƌ�&����˨+�1s<ǾC�	rU����k4�ʄ_�*KCQ����R���X�:�������=O�z?�G�(��A�Ço�mU��s/����Xt��Q-��w��~��W������ؠ�W�B�?��$fI��M羈�/b�,K�<qǩ�%=Fi8	lFAC��(x#�U�r[@k !���4������aVYl����~��ɂ=���Fl�J@�� Ћ�ᦗҊ"7�T0���U�o�U���P�����F~f��E(�'��{�`�a�Os���5�\h'�����I�̒n�~s�h����Zd�^U��#���H^�g6�T'U���Pqha�jl���g ��*T�T0J5x~>k.#�s�,R٠�zہ��ҙ�sf�;��i"$�u�F�h)M5�+�H@m428�Uk��ױ4,]��T��.]��4i�IC[�
�ԅz��iV�Zyժu6w����a=�oV�㢨�b��i'�p�}��ni8f�[�n�W��ǌH�C�� 6�(���zȸ(�y��FY"�W�yV�=����svS��*gUtQ;&�� �JJ�8��l2R�n(d�ߧ�G�}������^k]~��s��7�qBV;W�M`�*X���3a �	#� knN�f����ꫯ�ǚ��]�kJJ`T��=Gu=�Fi۶��t�IM&$�|��=�������s�/m`�KAQ-��]T���
	��lvņf2M�A0$
�N Ւ{��}ِ��-'�9P�j�~"-�R�))l�K�H��5l��`?0f,Nl�}a�ڲ�
A48�ƽ'��LL�}�@-	���31�.^g�z�'��0��a��=R�q������\���d���ߪQ"B&��87�� X+�WXL��3{{�t_��Q�㛫�T%l$@�}	l�[�-�p!�S���G�m�:HF���N>�H�SQVά�԰Y�5]��n ���R�p,�߭��Ϡ:�,/B���5�����vJ9_q�P3��
X���������	��z�X�g��S�V�ߨ1�7�����Q�U�Yd�&`iH�ڮ]{�����YЦ���X]իb�s��L��q�{�}XA�5!祣��~*xs�x�k���DO�U��U��u�Y��{±�=���3���q�٦�#���$���H8x:utjO;ʯ��gE�4�����`-�� ��r[�؈SO��]��֝��0�N�j[�t��y�qv�0;`��쾇�@�?�tnN����8��} �c|��k~�B���k�E�߫X�٩�IG���Us����]tIS�*V�k~V�|���6��Bso����<;�c��{�z�~2U�Sl6��bM�cZT��m$t����U_#D���ʓk��,Ҥtv��s�v�mi7��f&���0a��I �PEF��^�0#�	���B���P��������o�kY�}}R�J��Ȝ<�KY�ۥ��|�v�!C\ɬ
R����[��Cc|MQx7/#=����|Vͦ�@��O��}?n��Zbn��٬�J˒�@S���R��H�=.)���ܪ�|��d{��i܆W�3y��
�(���9rzz}��Ul>�XgU5����~�:�h���Crl������c��a�MG��BW��T}Q��Pz����4���ܟ  wU�� X%�m�*V�X��S_��1�A� @�R}��n�4��q<]$u�ҕ8�M �9�-	:���4�ubs*8VU��Ln�
�5��#G�����8���+�����ڽ��v���ci�Cf�u �6���F�%9��n��(\�p�x��d
 y~���g7�i~���yd,)4Dщ��CT u��n`{�hw��+��B���	3�m~�*X��d��j�,�d���!���ߊ���n�x����?��S�u�P�z�?qU�n�|�W�H�쨣��kL_S�u��Ϡ
o���Ҷ����H�*!��v����ߩ��IH#q
0����-5E����/�������lٚR2H5򢑋@���k�|�}t]ƃ�?��d�v���O�F���0�pb�`|�5�V�Sj�D��������T�#�=��l�#+^�1�q�d������N�������5HA��=.aD�-��7&}j+K�S2��@Ū�>�_S�*FN�x8	�� �OE��3�	W�1Ꮹ�`7_w��O�y�������QP89�F��if?� 6�NF��xO�^���o:�h�9❱��aU{x�%���X{8
�����Z��S��P�+���7ǉ ��Xի����j70n�6` z�j7�?��So�Ǫ���m�6:��@5��`-��v�xI�㢹e��'�,�����ߚc��q�m��N;�<�@[�r�K��k8��mX���]�vu*X�7��K�<�^	������-��<7VNTJˊ<wU��tj]�v�Eg۠�����-%�5=�T��]l�g�/�k�N�DRE�A�l
4]1i���c{�UTp4�f�.w*X��:7�.��
k߮�S�_|�S�qn�M���@�Zb��#`UԠ��w��`�ۨ�*U�L�E����m������G��g$��C�W��A�6i��k���m3����^|����rͺC�|uh(Y�F��z�b#���p����\訊�A����\!xU�q�E9�y҂�+�oͱsO9ֆ�K�5]B$Y$���L-@%mᴖ�8�pA��=�v�*�K��"dx�hm�=5�-�xi*�rJF���Щ^��|�݁BB������,���&�X}-�}M�)�i:���k�O�A�
�T�n�㆐P��5���U��V�����lPT���'E~do{N��ۡ��r�G�K��c4�ϟ�lzj6,�i/�z���?Zkb׆�q�<�Sl�w�ο�(������H���QoX���,�N��O?݁U�*`]�|��涮�����T�P��q�_�L2�W�'XZ'*V�5+)�~���I�Byg��vr���Gۊ�k� [Z4�������k/�8��>��疖��jԹ�>v����W[_TɼT'4@7���/�m�Z�X%^��FJ�JI�V�ۜ{���cm�bS��Ys�
�gW���>n�$�
{�2�P��[�:��)�w!|�j	���:�t��`�v�
���ʰ��S��X0+�@����~v��e������{������[4]}�tzs�U�ŉ"��;&�Ix��ڨ�pf+hk�/ꡚ��+�Rc\��*���j���~�!-�,b${w�vӈz�n�҃8�lh�c4g*Z��u��Y����`�umc�Q�@wj��4����2�P1E.�}������ٲ�-�e[�{:?�� �����:2�0�
eO� `�hM�h
�i��{��pWU�ה��zw�\cLJ��em��C��X G�Z��7��3�$��
$)�U�W�H׊�U����mm���o<�\`i(��=��ׯ_k�[���?N*l��o�c�~}�:��3[�v�U"�K����X-���!�5V�́�;-����mTpX�
Xe#�?�M
��C�~�Ӄα���T���8`�b-��F�zȁC �<�X\`�s��K�������&��S�`7� ��Rݵmgw�����Fw$�?��{����ٗ_�L��^�ɬ�F(5#��X�]iwM��c�D��*�4������~���k�/	y��5�����
�]	�Œ�zKMja6�T(��Am��z���X5v�+6n;po'��6�,��xʒ�d]Z������n���/_}{����G-.��5��(�!p���P)c/ꍊ&��`J	*��ZU�!
fGY�.���Q�+K�b�(��f�l�q� 0Ⱥ�i�||@��>�-"�#+d!~g�{�é��¥VB1�*;��ޛ1���pRk�y���|��k4 �ZUmDE�`]�=��x{{*�j�����cY	W5�s�,}<1�X��C6N�5H�����ͳ�L��ߔx��έ�Y���rmR��b5�)���V���S���sc�r���*e�2�TG�5��M5J��8��F7��^�Ǌ*X�%Y�x���{�o!�\̀$�V)�5�Z^B}����?8��bU��`%
���l�9�U�ھ�ʍ5oAXI�@Ś�uO����d5�]��u��/���?����_�M�]��B;h�`���cm���y��W^{��o��������J��EQG�����W��L�[���O�T�qi�:�PWF�!�ʄ_=VU�Y ����f~��e��S~�F"ZTT}��{ٲeM�e�f�)(6.T���fW���y�x�0��0�'4As����&�~���s���5���/��9�Le��b��E H4�f>˹���J���|�Z���������3�U�X��k�|�Hl.���Z\��0���l�Z�Kהؓ��m��Yd�чĥd0O��/�P��Y�[7;���l`�l�Qz����v���c�J��;z���6�Wl-��a&*'���Q ��(Nm.���o���mVU`�{���C|� �^�Yz(߫s5G�6V
wJ�<�i��h%`�J5��^ƽ,�>��xmp�g�1ʬ\��I�2��f��Ҥ����:M&����yIy�m��	�[o�|�o��Y�@P�*'Q�z֍WCQ�Ҿ����	�W>������܌
���g�i��S�́U�+�e��kh��?�Ӯ}R�h�_��:�`����-�� �K�^�Ŕ���.0�y�����x�I�x��go����Bl�R�1�t���6��>dW�p�b�P� w�뺎��Q��l�c{�U=V5��h�<�F�KJ���N��8nj9/e���χ=V7�֜�O�]T��1�y{����!Z�X�[MZ��-6��[�R��/W�`jD#*_6�p�,Ę��?\�1�ɇ���Ȭ��r6�LpkD�����
����|�E[�l��\yU������uH��`����UI,C��3�m{dyF��1�Kb�OcAe�a6�Q+�Az��/��	�آU�X�@�L��5k�)��?o\�!a=|���x �[k�-�f�B�N�EF]T��K�!����~�%���L�m���P�i%�޿,���½)��fy��K��ڲ)O6TMo�3�пq5V�Ε�	N����o�M"ࣣ���������Ϝ��T9�Z�۽��nC�; ��0-���M|�m�*|r1�����
X�;�x���S��k�c����H� �ty����-��Z�+�V�v*X���\
:<���>��ڮ�k]*�7�\5�aa�E�m��U�:�U���Z�zup�6�c�Lr��ؾ���<T|!������У�u�����
֭�q#��ﾻ�:�X�2c�=��x� ��P�!j�Y�#O��WYfn{��ݣ��� �%L���D������
�"��XC�`kZ�W�Xq2QŪ��dE�ġ����^K�5�>�f��kK��pɄ�69�U��
{��T�?^p�B�@��G�U٘ܖ�T�rF(zu̳��i};fYK
���П@I^|Q��9U�r����=i�,q0�Y�on>=�K�2�	p�~<�}�$>�z�
Jr2R���M��<k�x�Y�Km�K�Ù0s@`#�qU�����<�Խl�5v��WOf�Quk�Ҏ?d?;����ȭ&��Xͨש�RV#*�����s?�B��i�ڻCb�4�꫰ �]���� V��'+:0�����.��߸�TE
@��IZ�+U�sd�F�Xջ�/�P)1�4u$��'�`�>8�N��"[���h�\�g/[�<�F?�"N|llT��d;�� �ы�]��f���5�:Ȧbu��JX�X�4�M��+X�ڔn�&2Ǻ���[-:�-kj���{�\Ϻ7�k �fM��4ns�g8�f�{��-�]eXe4U���@�S�N����-X���	��
���o)�@��կ��8�8k��- :uH�;{�=��K�N�EN;R�/�~�M��+.8����ƿ������a_��J�ڃ�+�:����$I�!u�(�&xl�y滚=ж��g����$�]h�f��f�������j����5k���� �662�P��"��$/k�K�{+7 �hժ���}���8
4�?هo�a\�	�������4@N��K�y=}ܦ������G]SR�M�%�:-Y)4�ѽU;�������VY8�m�F�!W�6���Xq����t�Ͽ��H��b��%��3�3�sxg�r��p��֞uEģ*-O�bW��/|'��O��ؗ߶���,6m����F�q�{�3bLo�P�xQ�(�S�l{��ã��k*]������=�4捼���?'��]+m`v�ʸ
�M�B`��cw*��"c��� 6�{W��>v��G���� V�ף?���Ԝ
v�J����R#a�Zy���u����ğ>���m��٤�<���e���'��K�ۘg?��o�o�JhMx���ѓu`�b��RU�S�
:�գ��X�qt6�M���)^
>pLDԴG_�PaE�x�3�B �AM�t���V`�jX֍���u[�U>QA���L{w�U�g���A�
^�~}S��n����X�!��W��Z�h)�1�l���R�h:�X��W�����j�1x�7l9j<�P����iv41�(�Gp�7v˄��-n<}5��X.p�F��EY�V����? Z]�
F�W"�͹����Ɔ�%�u���
ե.�$@TsP���Y�������2S�X�|��تue�� � �� %l�oE˿��zv��b�-����S�9���+8F�sy��~�]3>��1�ϵk�}3�G�kp�كy�U�6���B���κ�����`�� '��蛢������}� ��?Z�X�l�묊�8�H�{��?D��du
Sb�E(Ϋ��WUGX�n��+��fK�N0���
�,JE���U�egk�;�p,t�*��K׈��@�W��܊Ͽ6�^|�]h`ăгU�։�uB���хܢ<+j��E����ː�P�����-�q��6ǎ;|��x�~�>�k�x�h��Lb�P����o/L�i�=��U!�KCcQk5��X�"���б�!U0�T��X�iK[t3��\0�e�媙OmP�sZz���s�´g_�mN���~�>�4��gdyǟ�d��5����F���YY8���:�;ЙT�aJ*8UpFj�]�ܳ����G��
.�^�T�d����F�S�N*�u�u�km%��*7 VU�Fǩ�	�ڳ��e�`�����q)�?�X��jX(�:���˶j94rr��{����Թ���O'��-F<=�1s�^�f��&�"1C��1'O6��A�H'p`B)�.GsV�qe�D���1�Q%�� ճ�u�3Iك�(i����.���>��[C���jF������RWG;�*nzݔZ���I5��b���f�p�U�qV���Ӱ��`I�5F$����.�:��II�\t]i�U�F$tne��"%��U=Vy�
�������]���k���Uƽ�Yr���$��z�q\��pa��H��Fb�t�Tp?h�um�Z�:U�"}�~��F�6���R;����CG�DM��i 5��#�څ'lm1�-˖�����e��~��E̚�i�?�mx'�$#_#$��w�h)�P�(J�5!�깒�S���7���u�:~�ƨ�2�D>����iP�{�i�ղv�� B,�o>#9O����QE'd�����S��v �Ƌ��!`�G<�
�P��eP�=�t"�*+d�Sg�%�k0��-���(������n��fW_s1b�z{����5��{��a^x���Xa�%�5�)���P�P_���Q:����'<�FT��W\�A�!,�cs�MLd�`�'ݺ���mq��(clj�̝PK�4�j�2���= V�����8XP�a���jOk�l��
儣JRբ�_��,�ao�y�5|S2z��X��qx�u�a'YF��VJ5�8'1ly��j�9�bB�/崪ٙ���e�VL�{��"�LK݋x    IDATJ�wSıH�ƪV �5�5��Mӈ�[/�=�>W=
5�㸁��U>l%`�(E�Rs��)�7㗪���H�!�z�גj��-�Xח8��T�DVQ�J��jܦC�N�.^���uy���$c<�A�^?Ѷ�J=	3v�X��,�P%�,ށU�q��D����es���֔8_+�ΨJ��LH�S��/�)�q�ۑΞM6=�2���HS�D����kj
����v��a�FX>!�!V�je�ŧe�=�xZ>�M��@=�����î��L�����6&Q�b�t���b��k6oE>#0i�N�X�f�,ST@#���*Q�O�Đz�T1��k h�YE󺽪�6���6>g�4eX7vhe�8��L"�{�S�H"*x���[B��1�ۻ��2M4�z^g�����:��MJ�����Km�bZ�O������=�XD�%n�ӿ�g���������8�N~���6�&c�bп�}:s�����+��"�h����y<��9��۬�� `@��k��m<ݦ-Λ����k�2l�}W�Uz�^}-�x�J���_��} �j/��NV�ZҢ#�	X��c��Hժ�V�a��D�E�Ӱ��r�Lf�S���ߦ����kIw���Q�(�?��T�o%a���ڨ\CY��V��#��'k�[���`3AqK<U�M[�횹��oK��@oN;UQ�p'��|be���a1H��7u��j٩��I7-\��O��3��������MRu!��k֍�>N�l�k��qD�u����yi�O��c�#YV��\�_�	�`�t���9����Oz�^y�u�T�*6.
���~L�.祝���
���aVu�?�����ꋣ¹�r 0Ǿ�z�=��8@M�/�M��S�]T�z��l#Fk@�ۿ?j��[e�9m}T���l�՘j�]Q�fa��Qځ�8� f�f�R;�[�L^܎o����Y[Q��Lj���Ve
/�/롄M2� ˆ����������C��PE�Ag�zQ�������=����h��-�����i��I�p��jU�9��u��/�_���-����$�W�-�/�ϫj-e�E��N���x
x�������N8�8���\E�'�|���WM��#�(�>q2v۴̲5�Q�S��x�e��SoٻdO+BOk4����!Ѣ��'�q�>)�F���SA�֖*VY�v�������R/*�1]�����vNź%`2�+Ӧ�>�l���ntY0et I��b2��^�ۨ�ZJU�7��*j�s2jd?��D���k��IF�y�:Yk��y�h�
��5��oT)~�WO�nտV��
�`���M �C	ZkmZeX^Kl$|Y*Ơ�/���U�B2U�"��Tْ5�욹!%�r��@bu��t������ �L�ՐW�b�q�b�Uy�5.��r7�<k�,��At��Xe��S/��:�vz@��04�>c����&�79/��q��ۥ
�V��a~ϕ�ܯR]�'Pp ������d�4���/s��YW�VT�����c���*��X�L�~�{쓅�-1����t��R5&BW����?̮<�KQ��A��ϰ$��Xkw=�8!��8K�T�y�������\<%.�S�0F˿���cxZC���YO� ݈*cў�rbdF�̢�+�mv��x鹶O�v�e&>��*�a1qE��W?��^y�k=���A`�v k0n�m����6�����Ӧ!���R�+T��{��ǋ1q��Uz��<�F�y�*J��J��lҼ.'�����FOáK`��CJ��H�	 W�]d3_��L�/��\
�����>�E>�wU����ٽ��i��+VQ���!���i�*U�wQ�]�v���݁D&A�x���BJ<6G{�E �_�O�*_Hɵ�:�R��A�Y��<�1��$�n�����^�� Q�P��(�\?�^��f�4��99.�j��z��R�9��=�*T7��4�X���'*�n'=� ��m��	�M��$c|�/����|����q��܍�u����5�|������M��&`�*8�cm`H�-}��e�3�9V��Lf'�d8n�SV];aL�*�Ν;{L�έ�q�?x��XS����IB��ڦ�W�J��%^ڶE��-�j02"'1��H�}��
-^c��q��w���5$���3\�I�r㩰�[���}�0�R�:�RUni@�V���i���/���PC����%.+��
��p�C6�p�����Ѝa�&��Z@}�$A̗��xFn\)�:һGg��1�U%�bu�JFr":�X�
��x�9�����.�*�D�Ԣ�K�׶�ۛ��n-�hkӁvC�Fb�kxs���o�z��& >;��K���'Eշ�$X��L&�Rkf"8�#k����;*�]bL�� f����`�g�zv ��E�X[���*U���V�"`u7%6Q!��
��*^�u%��g:��b���Y��O����T�¬.��[K�]�̪X+���j:�̝S���6�SK�$U�z�_��;������y�Q Cp�ͣ�=��������l��X�[۠aéX�Z7�̲E��˨��ZK�^�E�o�I�@Z���i�+H����^�z�e�^5`#kC��Ļ� �O@H���fJ ����e'VC������:��>*���n
�F{W+�~�L]L1��N�<��|{�����C��7�������h�`2CcXXT��^�Rײco���.��R�
V�U���&O	ܞ�	����I?B!��]_r�:��#}ä��?�^�y��l����5n�֮����!��Z8w��=�����+���;�k|����k���r�c�+}�)G��}�&3�:�M3��;DtD|%jNy�jS���`�]p�v����X#���|@ ��9?<��d{��eۮV�=����M!f-\o�JPa��M�dT�(n<���F�o�"_��z���m�3��	ێj\��^X�Xsj��|>_�`Z$v�!ôuv�._�v���<�r�7 `E�E�E��(���>�g�����	��αn��:�_�w�[�ڮ����}��rm]pH\��t�C�S/]��ivܑ�ZA�%��h�<)G��J`�6ƕJ1�{S���M���K���Rv�,/��vݺ5ޗwV+�-�v�����#�Z�r��_���gI ���w�x�w�R�mf��sα}���>��S?(�����E��ct�U��\Ԓc�b]�|��"��p^:�4K��ߊ=z	 ը������4��J������dyW�Z�+��_�'����"���{�P�n��ږ�NB�F\V��q6ґs��X�D>5%�U��r��rN$;��F�f=����/��?���w�:�^yo	v� �gNUǏ�t4��b<��1V!q�ϱ*6N&�W�!�j��嗏���L��c���^�O�bSDt��uIb9Q�����>���}Ω`�X���qk,7�.*x��͝�����ɩ"%�

��R�I/�uBL�����}#��~���􍹼����<`o�R��k��??b���/�~ё3h�E�6�mW�c��k�4k2�'6IY&z�^��~���1d��D�[�ȋ���c��*T�U�R�J�A�̲��Qd��p�ܗ��k�k���^�
�6.�GU���R���#�s�k�F�D�d��Ϸ^c:�Z
W�%�,����`�����O��*�W4i��5�c�u�N4���ZSU��G1�2�H8���H��������!�ͪ_�"�>�~?d��p����>����UE����u��x�9���`���Q��r����{����m�:&�[�|	}����?���So��O�~��R7i�?n9r�"��$�3&����<�<�cc��gh�������n]�Z��V�;��x�e̱��Y�#��n�;=VU��:ء�pr|��Y�^�,�ݑ�{2�VRRb�̷2v���t@{w�袤e+��z��p,�ӟ�ԡ�m(*�b��m[a��Z�����j�5�M�lXOo�����+���l]*�n����-��y��Бo���k.��O<�^����~�)_�c���X��Xo��F[��B'�����+X&����o�k�\r��z�_}��S�2�"~�y�>��y�ŗ��<V}M7���Mu*X�*��*VD� ���۵f��_M+m�(��46��n�/��46�G������f�C<��x�r�_h�.�y�2~^��zL"���J9w�K�^��X&������8HѪ�2t�__�uʀ�Q�L <�F�1����'b�@_W")[QԚW�:��>�q��MA�X͆;��z�0`��͗�A�����=?q��{̋��ՙ�~Ph8��	��!��b]m�8�Y
��[}I��~��v�هZ��Ѓ�J�am�d�`-E�w?e�<��E0�Lv�~�-�b���轛���?�X����A�Ia�[�	�?���%�.�o=G`�<��,���G��x��K;���O�YdMq4r=ĢtҘb�F��1N���*&؀(e�6��6�fƹ�;�f��M8���P�!u���s��O%݆d$�s�ե�|c�F�C��G��Xw4��1�)�UJ�XCʷyo�~$�A��j� \�(�6 �I���f�:)T���L�w��6�=���c{�1��,����Ʒm»�l�}��+/<z���OVٽ?��P4�{v�`�s�}��'����P�v�)'�q�t��k �zz&P0�\+��6����ΤlՆR��kc�ub�>^s�H;j�ζfY�=��˾+����۽�O�qؑ5��,X�[/�����c��5��t��XE+�\y�����J�$vC��F+?����]�**xذa��fd���l���|����L�3P��*
�)or�A���ɭ~~7�Tle�fcd�"� Z&�a�e����ԍ!j�b�L�~b��N��;o�N��{�*)���.OH��lu�J;�=톋N�́7`���z���=��2���wC�%�]$�&�S���Z�� ���`��RK���^e��ɏã/�m�M+��d�xkI��Ϥd��3hDG���{��թp���� �}�u���-�%����*��<���6�3w�k���h9lJ�L������޼��G��	��z�͂?"��m-���6���'���62���ֲѨAm�P�e׏Ek
@\S�¾x�1<��8<T��H�-&�[�xJ"�-Q��1v��ZI�?�I�:wJ��Xw;|��X�t�����O�vTźh�b��q�N�be�Ue�l�Q�V#����l�=z���o�O���rN�VP��ՙL*d�=�I6`��m��+�M�h�����{�C��6x@_���#����{��F0�.��ܿ�������EM��/�e��֧�?z�-]$|���Z��Uء���[�?�Z����e"�����y�%{z8SNI��`?ɸN��.^R�5a�ve�X�/	X%^|�E�X^n������wpV����S�zzS@PD�"��NPl�aW4���FK�bC,��ذ"Xb)�{g�����}�.X���x��0s��)���.k�%`��Ŧ��{��s�"AHsذa�ژ��$+��V�z�E����C^��g��}�Fn�̨�2w��%QZ�rzb�-M�XxnX.�l�Sa����M*
V�Q%�:��t}>�Le`����F�GD`�)#�������D�J�j�M�E|��m~n��T����� {PmE�uh��2Sa���P�U�#�^*�y��c����z��ڤ��y�����c�g�)V��^�,�u��k	���,�8�-j�P~�9MS�7cϵ���%V��^�H2���D�u�o��MO��m�a��}�U��4"�3V�Ϩ��ɞ!�6����RŒJo��t��e������*�W�(E�=V%4	j+R�L$*R���?&�@��<�rR	Zɤ>�*2w�#IC_%z�"��9r����DH���W2��R�>��mܶ7�#5�=�2��ɡ��ցuѲŶ�/�n�Ѿ3e��@lگO/��D{��Y6�)DH%eG�m-[}]m���(W�X�]��+N�g�xO���н宇�#^f}��嗞c'~h�?��!�ջg;��/�٪|BfPU����y؀>v�#��7f��/�f���C�/-Ɲ)�c�����7��!Y�ǯ������W��dA����F���J��0�*�����$i(��m4�*��m��f8+�5�HF�ӧO�O?��"4'����ۄkF���q�#FxJ�J�Ͽ�23�<I�Y[������߅Ν�vWg��W��@�G8@�(�9�6�-��Ѷ*�z�\u��J�&�e}uds�E���㟲�KQq��1CE�&kļ���a�Љ 6h�k$^C	5��٬���{��u ��*�0����O����=�d���.N����ޠSm?��7��1��ͱɶ��̧�Eꢺ=VtL�{�a�>���@����ȿ|i5rHU,	B�﮹����+�G1*��%�g�����᧭<�9O�b�t����,`���;#��q�YL&�R(�*{v+��N^�f�!��zh������G#�0u���$W��hnW�|���/�`몂�6]=V�XY-i���S�U�,��S���=$"��Ey)8�p� ^�n� ;WR"? X%����pI���)¿��O~����]n�%*El��S���U~��S
����5v�y�ځ�{ڝ#�\��#JO4�3�+��n,���#�b6UZ/�27\u��s�T8�=�G�ǃv�=�b���.��<{{�d{��w���\��[�Vv�_�rW�x�:�ҍ�,���5=��o��aQWB�  �$c0Xo�P��M6Ny�m#c8u���ѧ�`�";񐓒��Gyi�bW^�:�?�R^
��3Ғm��QU�f���"̔�y�h��������eKZ���_�9�`��/�R�3�ew7:/Q_��fϸͮ�A)8���S)�����<+��O�����*-"�~�F���R`���^�[[6������[��&���3���եgۑ���}|�c�t죯���}����*D&��05B*`s�(;x������x,Yg6sx<�a�^%E�]Vy��[� R��e�|8۞|�����)�����FW������M(1 �N<��]۵�"t�Sf��?�7�6�q��?��K?X�kY6a��֞+����,3Ռd�~o����bS�s����z�DX���[��>f+�*�q5����XI�5e�����ܵ�,�M0&$q;����j��#�`)/�r��-����>���wḼ�=��^��]�hw���ȑ#z���+sG�ζ�ڶu;�'5[2����۸t2�2�0-��F���Po��/�lֲU�2�MKء�g~)�e�b�r�|�M���.�u��ϴ�^x�癎?�d}������%즛�'˙hN��AvC}��l��>������55=�|˨ȷ_BhA9��~m��?�c�r��ݭ�w�Z7���b�.�y8#�0��I����qqEf�
N�^o�	X�6C^z�b��%��V�l�$�_�j��&c&��MQ���4���7�[2���\ł؝_�"���<YM3j�R��
����l��ٝ-�ވ�UZ�{��w�ա�E�	7YP ����H����ɪ�8%!�g��K7o��[aml雃~62v�:�`��ho��#x�2a@�R>t��C.����m��98�3�2-�� �gS���[�{cy�P�Q�s��q��XO�d�̴����q�&Ӂ��O>�������Sf�+��#�����z%�&��g�!��27�xd�����6p��D~Ip���6��7i��?�I�V��㞴"~s-�����H��]=V݃�hD4(�E���*�^�M9��+.�'��R��9/���D�'Gd����Q�Ӭ�Z�z������:.S���/`��֓� �`P��n��5~.�~��-E�833�q�C���`���P^�V��ofa�@�.I�)cu`���wr���W�u{�rx3��+�\������� Xˉl{/X    IDAT+1
>�������y�����Ղc�>��[؉G���_�b�`%�߁v���e���L�ؙq�n������oy��7�s{�͉��y�Y���=:��),YO���
�SZ&�ڝ���[CD��۬�~��I'�d}:g"���T�RyF�|ޢB{��O�-��k�ג�)��6IU ���X�
��M3�*X������\��ZTU,������F�q�'(c��E�}�P��
P�/_�`�rOT	�b��lZ�m���R~��z�N���fW�Xm�b�Q���A�vF(�gE&k�44����x� �C�5=���{~R�:s!�O�h+x�$�h�SuJ.]kW�{���q�>�˪jKAҳ;ky���v��B�QL H�^�U��K�e6z�2� 䫔�"�W	2����r;�O���ƽ�O{���4n�L"h��IX�����8B��s�\�y������+�#co��<d��2
ޜ<����q��������4���h}D���.��!a��i�_V��:ѱ]J���F^A����ྴM��������UAOu�J����l���Ͳ��c�L]�ۋ/��x�F'w�:}VL՛ B �2�*܋�����K�?X��
�^)8��nE^Bd^�Z �D�d���X��� c�w��m��u?��6l��;G�E�*A@(-�h�����|{g�?m�Ï�AF6�t��ޱ>�ӏ�.K�k�^�3�ڠ���o��o�u��ww�=n
�֢���Ҋ�!˒~������m�?���*��n����MAf��V�a��jRrnӆ�"�����'���+�bʵ�幊�x"�5��VX�ŧ�S���SQk�rU���YJ����Ŏ���6Z�;���Wf�A٫�TU����z��J�"/��b������;m�A��ƥe���EFn(�C���PUR��Y,*��C�>5R�R����ϵ��|a�ϘϾ � 8�1<{֘�ev�Y���G��l�Ϡ*�)7��M�v���ی%��Ҵ�`)A�5A�QvT�j�Rs��2�f������K�e���M?�6/�|��ε{ �@�Vr���^����	L�	��YE=X�<�(/Xg{wȶ�_{��4��-�O%�-���oO�qϼf5i�=x�&��^$c��Ҧ�U����*��2T���s2�ɼJb1�ؼ�n�3n2����j]7�����͎V��Ha�\�*v���K��g���G!˽Rߛ�H�2�y��G�P	dL����Q�OJ�>n#`}�)�iѢ��:z\�6w�l{�1����Fl�I�z��-z�荦q'����Â��{3����2����nS���fܦur�Go�}��X���X=����6s�I.�z�6p�@7:׸�ڵ�xi��Ë��~�f�(������ŋ-_s�̐2����J����B�ߧ;��aֈ��������\S�yK`��ݷ��dH7ʾ��k/�b�`�_�=��[���_�ۙAۦ��o7\v��g���<K5劋�@�ogoc(��F��:��AkC�^z�u����l����LQP7d��6S�x�
"Pi,h ���F2k�b�N�c�?��$�܄8-~�����D�K�&<�d�X�*K+XF�i��Ws�rǉ'�
��)ٺ�|���>n�3��)�6����5$Q�Df�6C!�`�"�mo��+���6ߓ��0뒆��_#[I�lVQκ�Ԙ�v�FH)���&��@J�G �w�.��l� YS���?����q��h�$�j�=��E(���#gx���sN�,�����d��/s>��������n��qi�{�Z�Jzk�Z�r��Q��J�	T������m@�tw�y����3/Q�nn����gD�Ȣ2�u��%����A/���Q�v��l�����cQ`%,�{�ޚ�է!�}R���q̱^3�R���O����5*� ��~b�f�6z�P�Fկ�@,e5��dF?�
i?�m�q�y�b�6���E Y�]?e��~E�p$����h�c���G?u�EcH����o�T�m�O��Ӈۄ>�7ߛ��W>��9�]�=�L�Ky�b�c�����)3��Z��mQ����m�R�Q��ч��"�z���~�5��,J�U>$��?2[=|֜x2��� B�T�Y��Cb�)��6��w�*bm�, I��U(�����p�g_|�Z���K:�h�����q1����"[�b%B���2?�ϑ'Y��,�'-���Hos �ճSG�#�Nܠ%kV��?�r��^g��vf��@��/��9��)i~q~�e�8w� �r��/��$FW�S����� �Jz�	�{W��]�`*>�+�[�E���^f��`������߉l9�Q_c�̱��<��=k�}0-��r���'ҬZ)-���I��X/sV�8W^
�m��
�55{8��0+�r��K
DZ�[�N�KZ��;yI����Rj[ll�X�P�
U�B?�"�*�*r��C|]�K{�mvE8�rLV��:���~ �
�&)֮y�?d��3�ǈ���W3��w�HL�r����$6�D6�J6>��!2֩o�}`�Ye�Z�۩������2aH&]�m&�g|�ӹ����aIM[���+%^ �_%^bKh#���ʞ��%ˑ,��K(��g��c|���4Vw�!�efVUP0�𜓒;�j�KD�<Vd;��� Z]��lh��&�&'x�%����(���u�_����Y|z3��|�Ƥ#\	4C �BA�cV���z���g���P��ʑ��]��j���4�V����N��*�z�
�=��A���J�Tf����w�A���.����C0r(U��޺�ki��o�|m�0�!��z�s�.�D(�M�6�n3��yd��6�s���UF���$I�Ԫpv+p���={�"�һ��+�V,�u����)�
�󔮳�=ꕻd�Vg~i�h'�:x�`Go��U�/�1���M�P�U�QƱh���(���t0>�e����ˢ#�s���v�b�(�6n�bMТ��3���c+�4�ȢK�x%-I���q#Kx�a'��e���|bx����{�>]��>ir&���1J��,цg�!�vƩ��iG��O�Zf���N�%��J��^��K8�v���`��mG5#y0b�����x	Dd���"4n#`�+��}��|-�fm<��-�KI B��Z�Ļ�K�'�Lӟ��%C�[��1C�qe���������X��'cݵWG��|�7@�rh<e�rRF�I���΋gmJ���n�is�����Y��k�%E&����
���YdYU�s�a&��T�s�T[l7^q�ܷ�e�����E��U�����Ӵfm�L�g�d�6��j6]q�k1W)���L���]!F�WI�xCa��V�P~� �<�b4J#c	8z*%h�ws�lpM�ذr�>��]�(k�V�]g���>kI1�y����EcV[���l����s�C�6d���z�P$(Ha�0%��ڋ�����i�r#Z�)�x�ŊƠ=擆�o�Мo���`�&��l���e����[�� X��r��l�$!�a��"g�#�zv�h�w6��M����5+����~�Ko�R��N�/`U��	�
� V�W�����Yݦ�֔2�1�Z�׼ys ���M��"��?uP���vNQ0Կ�ѫ�\?F��Kiͥ2����(g#$`E�MA�0M�h�|�_�X븈a)x�G�[�@O3�{������q�]��P�1T]
�g��ITi��>����X\F���Ĵ�meDr�sW̹T�To�!֠���#9�R`�J:,�WE�tvW#�#�W.�,�o&K;�����Z�e��,(�9&]p�9N�v��d��Rː���+�Fy���������̽�PA�A��y=���S{��ih���=V��֧,A�4"3 ���@�l��
N��+�^�D��M�6�d���X����kG����T����R�2V�hdt^Hp�Rpht�����w]p�=��N|��X�1�]Wb���ڿs����� �� g����eX��]�����-}�fΙoI�WEl �)�'w������N��R��RG�p��C
�������6􂉱� ?UJٌަ����0����߫ gm�.Ѯ� ��Ǿ!�f�W��,�o���c�����g�3(Gq)��-����n�AkH����`�j	s9�'^�dϾ���+I)=Y�A)8�0c��r��W�&v5����_�x�}��2K�n�F�aՈU�����z�5HHV��w���k1@�'�j�T�tϾ�^������I]Х�C��톼u��w��#�hDu��ɥm�'A*�!�Iho�S�k�Ry�0�U��QrE�U�m��w^���\�����1�Y'Z��̵	�Ū�A��< �J�&1�{���Y���f"[y�Q;�u�	V�����>W�_۽���8f�wZ
>����[_���X�*'�[�q��.�\FB�8gnE�5��{<K�d�:�pG7Z
��ot�����>����v}��p��z�^�Z������Q�;��|\My��Q.L�'��(Iw��xu���n�dP��y�^��\�u�ȋUH�%Y��*�C5X`�e��:3ޮ<s$e���0�����J�-�gv�~��-^gy�[���2R��I^
F���Ȯ�R��|'/%�50VE�%���ÊL'��޽'
S�^9�_3�������k�"׌6�i-�Ac�նl�*�H��ƅ=�Pyi�����c乬�H�ݒ��/��_ec��)m�z�<:���W,|.U"6F�[ [
�u�6�JX
ėzZ1ʬ$�W˿s�d���1�O�F'�}"��-���G%����ɘ�ZQY�\��JKeHU�\Ӗ
��	D�U.VA�˞�H�L�����%����Z)J��$T�#�� ���9�1T�F��Yr�r�Ay*��[���m����"K�6�F~�;VUx�y����fC�J�����l��y�W���޵�5�0GQU���SO�ܑ2��o��V� (��k\Iħh`�B
z��H�K҉�W���4!���(��BJ��/�:H�j�9��6x�a6e�{��7��Rkp�4�=V�v����k�e���v�i�Nk*o�֯6���G��
�*H�y��*�s՜�L�K��!���/�s��e�ߨŰX)݋����0;յ����� ���k�$&�������2m�Î����33��F0nQC�C�I���F��Ö8� ���
ʺL��4S	��R�J�*�4���:� t����%F+_ꤔV�r��O%��=��Y�H�!�S��d1�R��}}�L�J���������{�k�YF�.V�f�w�,��H)x�z���	��$��O�8w=Xr�	�γ��ۥ�^nͲ[4��|n%Ql�����6v�*����.I�#�����J��>���D�S=V��㛶qI�="�����Hj ?Q3�<�b��²�i��E�cټc�2!Y?@Mż8�<k����%�h>��U+\�A�Jx2R �)�)�=�.9�p�R^�n��UJK��#X����{����O������5���N:��A�U�d�L�9K�cT5L�3�QpȌ��E�ӗ�O�d�O��t�qC������]��� C%��F�|�3��[0S�LZ���sG���U�B��j�d���g�l#��[�r����Vz�Q�n��0a�:�ۇ_,���y�T3� �I�W���R�����bC%#��X��~s����G(�M��L~3jO�������,������
�oo���M��|����&M����� �"�H�5�*,-�������WM�|3g�7�z�pZ����`��L9]�B~/d��X�K����J��%�ƷQ�p��y(c���[�`P����*��&��v����L�s�HK�2��pH��9Ɂ���d*j�������Xt�zc���������X��0iFV�m-�.Hb<��yA��է�J���f}5��>'J�'�L��ZN��<y�EP�,̵t6�֭ZX��]Ț$��hkP�X�b��^� �RtN[v�f�聈��s�1��uW]f����ǟ�t��B�'p�VĈ��j�b���m�(W���~E�S�o��
m�w�M��_�JІ����Ώ;����4�� �<�B�5�95n�Gy��]����bN�'ʅ��U��욠��U#�FNR���� ~_C�%of�b�*��}���%�R�sZ*r��d�FU'Z>	2�]�2���Sc�G�Q���I�P<��h=(�����>�|՞Y[Id�"N	(���&�k>7�T�Fc8dݪ�US�vst�=�1�w�lx����=F�ŉXȍ���>�HkyRe��M��j�o��IU��|��Ԑ�6Q���S�� ~`+Xk �)�����h���ɮ��4됍99'�bE.AB	���U�l��ϥ]y�C�ڧ�WXr&u��5P��W�Qn�*�k_֨M�恕�`��W���y�uh�jO<���X��gj�o;��c �ͷ'�}��aK����$Eexe���X%iX+��w� �ܹs0K��sY�Ȅ�qۙ[�$ZG�ݺS!D̃�9V)1��l���ĸ�L��
� ��}g�u{�`1�B��V�6K��xTo�G��lyE>r�l^"���a/5�����W��E� '�H�g����H)mn�J�d�\P-z����Z��JY�I(`3sf���O) �V���K�!��M��s��D�.�,5%�i �2��N1 h�f̈��Xcxh��Zk��yKԻ��:��q�>�G	�e����g�ƈ�}��"�X�/)��ˮ��R[M�[���� �2�Џ5�k+`�γ���@�ܹX�d����hY翻�֔��H��.we���9���6.%-��U�ۦ]y��`�"j�����_����L
8%��q�BRu��H%$d�%���+؀�l������z�1�66�ڶ�f/Ze���:6���4'�%S�U3���|%�ϮR���EX��3FZ�f��g���/u�-�0H������>���-_�|բ�9��L�ڒ��i��GrT&UI�,I\�[���sα ���k��ig��8��YS��h�J�O����T%{�����>޾���-��R�KLa/��*�RX
�5��P������6��ٻ�����^�8�U����/��X��4��(�$x��v�!9M^�ʣD�I�c�]:ى#��2��6�9�	�SZ�1c�������"�Ջ��H��"�a�*o�M{�`gg�� k�ो�/���W�������*t�>b@ʆ�]��$N�;�9�P$��l���޼Q��$S������V)5�&��ڣ�;��]=��I
X�,�q��_~��z_!xz?��7[tt��hE�I ����`��C��a�Ү4��Ϡ�'>�,Lc1U�(�%W�Vpc�)�(�ʻb�j�����RN���a�D�˘�j��|�m����ג�@���Z
) I�K�7�3�9V�G��i2�T�d� Ѯ-�i�7��.ݭ.;ڪ���˙�z���4N#��Xgo@ �2[z�2���!��+�%i��X�`���6.��������i"�`��.���ZkN�U�G���?�l/�����
X�c+���R�e�Q^�>�_y��鱖E�9PΗ^�$;y^�K�a��S�_?��^��:0S��1�_���3ۻn�a�ÜO���i����E�'����B�:KL��ۮsjP�W;G�d�@<�����ڝ���^C��C�E�����/�����(u,�%,3
��Mm���<����k�1k?�Am�E��֯[';��c���s���l�!�:�|�F�~�c/3^4�v��dz86�B���2�0�Sƪq=	���'�/���}��֫#k�R�Z�l��\�,^�N��7n��O��*�w�kD�)�����f=��؝t�;d՛%ب%��3�,��䮶J�U��q򺍰�%��X��d�SF��cܦ�x=3��v����nl�7y�'���-�P#oj    IDAT5�Jl���g�"+�	şe˖�B�������t�f}�0�
O��M]�j����˛ ,�r�X5�*f��k֐�K��W���]���_oݺ�u�A[�]�@�Hg&��.R;���T)]p��(�j�K��(5��Y biU*�a��4,���Lad);�zn�nvU\]�-�5�9�2'*�}�DD*�Sb�<��rv���Lb����Z1O��$6����;����(l���0�#�.�f�Q~N�ǪR�*�����s�"6�~Fi=�c��MS�).��bV��h,i����`I���"����X���XM���������dS�}iϾ𢓗��չ��d�t�`ͱ����`����dڃElT/T$�#�=�Q���,�.���_�>��2�HJJl)H���ʦ�6D�̫�	/�nS �����ӎ���HIR�i��6�M�h4�25����c�Z��B�te^��`�H^��X��H��y�SgٴY�m-�oU��������*eq|f ��W�Ro�QC¡~q�6�֫{�گ��W+��8~ޛDP-v����ي�l`?y��-l�6W�2J�ְ�� ]@��;ǩ_�9���c�U�� "���m4������M� /�L�1"�����ޙͳ�m���xD�ֶ� \]�B{k�⤯S��������/���ɗ��H���
2�Z��Z�#�^�t&,���+m�+�S��	���g���?ej��hq4X�D�T介���"Ǧ"�2�93g��o�k���Jy)�X5�J������4�ɧ�ǀU��r�������ϯhx�tr�R���r^8�߾}V?m��-rIC� �2m/2ִ}�0%����PJ4��ۥE�KS�	�=��IzS�^��*�ʹ'����HҰ��dx?L?}=pK)����$� q�b���_���&��<p�r`�|�Av�IGZs���Jʪm!����[.vEy�w�6 0Qm+7��:��D��Y5�+6 !wz�O<�<��a�VpJ�RW^R�*`���K\���MW��޲V���a����{�x�F��
+!_|�O/˘�� %�� �m�
�X�!��� ��ĸ����:�4�2T ��-�5�-�t��~v�IC܀��<Sg/D��p��$PlKk``��0�5�o�hM�����ت�2�D�S%�*7�|�������)��R��k��Ç�	�[[�\Dz԰���)��)���v��-���Wق<�8^�&T��]�fc}�QKȒd��)_�jm];u��=:Z���r�U���j�F[�%��L���<�2.\�~D��j��Izޞ����Q"��@V�gq�%�ֶI*�c<���_ﰵ�i�q(���R(�j"�F'7���ovx>��)��􏣁5�� ����d5
�|�� � �Ǒd6 �"j�i~UA
�J�23�{��H��6����>ǅ�Ew9ֺRZV`�d)	x���
@$c�q�n
��H:������W��!��� .�w"{gB��`FkpW�	X����$c��A�`e��S�@%#�m��吭�n��ߣ�5��D�֏k*��rN.�T�1�:v�n�:�L1�{kއ�b�\��\[�|��n3G�e��?�d�k���M݁d�_�ֲ��Kc��!�z#=	��
"�<T���x�ΝokV��<��%c*ۈ��!v�ȡ�����	��NCVm�-[��g,7Qƨ�4T߸5��AE��'�'ĪD��X)#i�J�R^���U�6V��2x	D(hyƱ�mT
v&՝w�W4�\-e�Gy��/�>��c{��sM2���Fmz�k)�"����C\����W��yA@�FW��r2��/�έ3#��W��O�-ĸZ�5��L�j�Ӳ�]s��d��D�H�����:&	���ҭ�Ȉ\�I˥���a�a��>|	�t6��9��h]!�艊�N75f�<h<�*��S�W�#�%B>��m$�.(�s�1��>Wc�g���2BAJ<$�nu�2�@�Gx"�iYQ ӨB�"�@�}���ɗ��zkڢ;� ˥Y�G�u~���>8?��E���Rז���kϷ��ԩ��]F��L@��Ai���n���\�X��;m>��y�D��V���)��� �aL�5q*��R�U1�R�pj�>:F]U�1b1���L��(w�R^�����3d�:�F~� )���u�y�����I�Z2�T<c0�?`�iHfs]�YO�4�Rj�$�>��L��𝻯>���c=�S���R�(�*G�<U��ǢU���:t��5b���F�m2�$6�R�v�Cb�?�֭��JM���������ͳ��O=c�Q�8���s��u�1{���އ�����w�����|�{�v�*����X�'͡|D����ؕ����/�Xbo ԟ�JR<Xݻt����̂D��K;-pڌ���4���W\�\�%y6oE��2C�Dq�A,mBU���=�q���m$i(�%��X�8�cK��X�����g� D��6�́U�D%e�2.n׮�{��C�$��U�`	D��Ь�eR�Q)��{�z����vExu`��<�TU���A�X�a����n�~1��϶?��������A9W�
F��e�x��׮���d�z}�=��kÈLs-ω���ՆXG�1	�JШL�Ԕ�jX���g�Nġ��g�A��YU������/���1
<���=����_� @y@����b�~��EH\_�_���f����3�Zr:�*JڲQ󾡦�h����gi;���	�U{�H���[�4�q�9֯�$b��e���*�PX�,w����'}Faao&���c ��V� �胤!�*� 0Nm�
�5������T���
��5���V��`��x3�c���53譀�gYub�o V}���
"�������f�IC�����H�S�s��֓O>�9�/XW�\��u���3�`�����mq��{�߀�������XR�^�kڻc{�����W+���eT�~��H�x�2S���`a����Ge's�}���v ��:����z)�$ۿ_�����q��G�����\s�,�o��ŘB�[ӹ���a�3q��9k=�Чm�(W�X+�1f"bܺI#\(��O�ֳ� ���"���3�̵���JJC�IMo�f0G���5?���M�����mBICk��o2ֱc��HG�e����c��0 `�����I+��R�.]�Ǫ�+�y�_����N�Z~�)-r�7l�m�ôX��nW�S�ZKV-��ZؼRW�i)ݰ�ث�����,�L�7�����l�?Ԩ�.��l�<F)�:?���®��bC��&�9�y�=����O��i��˦2��L���b�&Ȗ������ a
�ďb��	Ϸ!}0dc5���KI)�P$�Ai5���\2OIS)3��h+L�":Iΐ�Ty�^��;�ޜ4�,�dL@$�)rT0���H�%"�XN�G��]�*V���p��PyI�/`��n��:����EW��ܧ;bi9�#HS��R�����z���E���JYZ@��kN�vƺ5����,�Z�i���
c8=*J�|M鹗G����2E���U]�g�����C�@�AY��DF����5$��SP�QR�z�e���� g�����G5�ӀC0R���艗�É��pu���?A^R�U��L��G��u��V�� ���i��/�bz�[J��Y2�6�X/?�l�����c�fX�m۶�}hpj�rRH�7R��n���Y����?�X��ow[G�0��n7�q�M�6�N~��w�0{�쓯�Z��-P��V-[a=��!������x�r;i�1v����G&��i3=R��/�P˂UܳSk��X�N9֥Wonn ��<%/�?۞Ɨ���z���;P��۸� �Fi��F���"/e����G�t��$i��e��5�
y��C)8Z`D����w����ٴ3��T�RWJ��
V���0{X��zw�/�������y�P
�O�V�v�؋�[�[O�}�Cl�?��0BAr1�TZ9u������}�X!�ރϽk�~0��5ە�ҥW�-�TI`���u2	���O9 ��|=Ѧ6������;�	{T�<������$%�t$]aRN\��������O��C�q�)��|MPQ��VؤOgػS��5p5�]ÜI2ղr)ɥ85���j�=�I��K(^����L��m�P^Rv	��Wάj;�T~��sa^V�c���/��97�=Y�H[:���/��L�ӽ��b�NԎ�V�������h�	C�ʹ�Ts���V]V��͉�N=��#T�܁�=��͖��79�م�\G]gL�l�\�R
�K�E��W��縒�W�1���gK!sI��B�.|��]�zuG���%��ۨ�6���E~}}��nwg���I�g~�.���7���cզ�ƅ������yV�<[�y�u�b[�R0i� �����AD?�~�˱�f�:���q����&����t�ҭ�K��@@R��t�F�8��Av�yG��o����]g��|��r��n�W/(N�Gǿ`|6�Z��p�//Ân���.%�)��}m�j�:�u8�|��"���m_��G9غ��,���2���|h��!;�'��R����6c�z�]�q�<��R�X��e���A$S�4�F��KP#���Z��ٰ�|ѨA^���4����f�|��������I=���F�`���o/��Z(�G`"r�Im�с�J��?O{2�]L��D�̈?��l"����������?ӆ�ۙ����'�NG����b��a�6-m�>=�b���,+��_�v�͇`��B���i=��	ؒ�J�M#0�UeY��vH}G���Be�"�����Y���� ������:�k� }0�)PTy4(���K�� �﹑S�F
�ߓ��r���Q	�z�fq�\�T��H�~i(ˈ�7�*{K�Qc�P�+�K�T3�;��6.X]\�r���T}�4˄u]o̳� ʿ:����1�����zug�!ݾ^�
� �YF�<����L���bx�
V����{<���AP�p��@؁�?]�N#K�F"����P5Y���ӹF����q�ą�5q_<��4<���j$�		�2L��N�V��2)�{�R6}�1�Z!k��ؒe���c@��b��
�뷁�T�5/��H����L'l�'���-�6�=��lȐ!h�����F��M/�.�υ}���j�h	XE^RT�l�R�+83���,]'Kk�̮��|_T����l�T�=v�+)���t��`�����:��C���G��{�>��cr�P��Q��ï�j��w7^a<������ֵC����������.�,}Eh���+�K��v�M���w��!�a;��3�QL>����=| ��a��h�{���H�P:�G��JMo�ۨ�_�P7Z�W�c]�WL)���N��+�zr1"�������6鯢9q�j�ͳ�Q��W��#Fd5�������^7�� q���#b���9VI���zI���ʫC���ɛ%Ύ�F˟����yЮ{1�IO5Vz�f���L&�W�H#8zV6����so�{��F��%��� ʔ�Ϫ/Z���`g��A(t��JZ�JjOl��r�v��g�.��J�����f��aq7�f#����^%�;��Kl5$�E���p^�4A��!uT�����E��E`Ŧ�f0���*�M����h�Q��FQ�3Q~�
D��*m_)/)��HMLD_B�V��
\K��l���3�PXXj���S�����-=k�3T��9`�AB"	���
��g��:�q�u����@Yef��T�w��{x�c�!VIL( � �C����Gl`�X52���xb��k��{#:�+�y�:�4_���m��J��X�X	�,��x+`=��Ѷ����p�z��6��p�4,�7�a��m/:���X��>-�.�"�e	�;Q"�d�"ݫ{K�˭��Z��E�D�w}�:yܡ������q<gڱ���m�=t���z�xƞy�iֳK7ڣ�q㟵�f/���8���+��ٝO�aqi�ָ	��k�u��9ݎ:� �띏���G�J�ւ�I���-_[hk�m=�	X�.[j��l\�"��ezPpŒ]��-��5׋��bʦ喿d�k�tFUF���ڄ�6��؁��h��7J����ЎP�F~�b��k>�F�j�D�2:Ol��{��k�4�'c�5�H���B|��Fq`�&���N��'k����b�%
ȴ�k\ ����¤|����v)_LUP�7���(p�f�2��G ʵb�E�����U�V��	����d#HЌ��U�4�	��u�-%�kmʫT	C�Z��Kn^��I���J���5�8I1�V22OfvNL��+T���F��EK
X%7��J%�6��2�:un*yb/uڊ9������I��֕I ����o�L\�臀i�)y �?���gP�����[��CnȄ���/t,���!i*B�ꊆ���y�������kY{����M��dj��v��
��,`��;��X3P�6��X��$J�?=y�4�u�ԩ��E�Hh��"��������ek׭w���2:��s_��gMs���8�t����P�H���h�.Y��2��h8�{��6x����;�n_~=ݎ?q��uڑv�����o�r5��.[�V��&~�$�w��}LϴM�,���3lͺ�v�8<0V)(�f�Ѓ���'d�MZ`�y�%Ѳ��wj�Vp�u���Zҟh�sm�����AgEJ���g�s�MD�����s�?��Ů���5�TJ`��WX�Y�����0��Ct�Rp˶X���G=���������5��%�8�)���5�@Z�����
N�nG��^��<�����	�q������3=D*�!�P�|hX��0�޻gw�Զ�ˍ���W��"f��ٗ�TW�QF�9�՚K��_D�>�qB`�lҍq��*ْE.W@҈��ʰ��2�S!J$"��V"K��L��9�	�K��Ȇ$Q(�Nٞg�*%�\#!T�!��3�� �mE�Ś�r,�PC`^]�ю:h�]8r����Ѧ���VTP��A#kپ	D1i���Ͼbo�s1��l�W���\�����C>��-�h���v�	�'�󗮳'�~�8fe*E%��_�����0�~;2����D7�\t2�[�G�T.��/��k��u����XŚ�
�:�惷�vط�mv�!33�Y�ߴ��Ӹ�)�e��oz��~��M@
P3�=�0cU4��*z��g}c��j(_�R��#�F�%P�J�O;���,��Ì��)��Lw_�}�jk�s�푧^���������~�Q�胯�7��X�&i�g�!�/<�g�w��:�a_XG����]`hM�G�S^�g����,&�5��[�l��S�!�tYaU�E^gO�����R�����E��eKJ)�!�����k�!����i����v2�DX�q�^	����F%+�h�7����\7U���2���V�de�k)C�ίp\+��F�y���7��U���!~��PҰ2�,6�=�]wu�V����K+�{�zV���Z�T0[.�*=���z���Id���~�:V�>�@�3�ZN@UK&%��j�J����Tj ���,6~�
6ހd��$�p}�CrjR9��ԥZ�^�`�j Fg�Fʖ �������<��� .�K>��KP�fC�.[Fg];�����@ĎK�;����M��\c��F��nMl��\{���}���s�t��G�~=��̕���[�[ae�ŦV��F��`�-,o�~#%]�c��9��� �Z	�e����U�g��/`Ԩ�7!,�z@��'�,�M�Iv�*רWf��н�� _��
�8bF(['׾�������*�T3_�X%d?��a�b;y�)�ɶ']Yd!P�ArOMFu>|�[�n�Yc����X�Pa)���*����֚��U�6e��]c+c�qF�+��1k�6��ޫ���r6�����S9C��������Ͽ�a!I�s�>=8���J�K��)M/FQ��ML�ed�t�\]���00�h-^��nH/��ΥIZ�5�鼱������Kkvw	g��s    IDATD�ǚo>+ao��J��k<=e��4$NK�8#ӁU�����%_e*��ܞ��돊���pf��c�@�$㚴n�c�C^ڵ�U��2k�A2qu"� /�D�/7�ՔV��*���Z�e���ꉩW�#<��j��D֨����݄�M4蕅��_�r��&=n}Y�tj}V.<
��бG�����!UIkT5D����@��z9O��b���}0��p3�n���k�ѹJ��@����� #����_�g��f���W���^�^}\}������l�O�%����	��m��%�̤B����ǿ��֠b��9�(PK�"�9�8��V����'�*���#E���"�i�F����AA_,{����H$f0Ɏ�7L��D��Rkޛx׵��K��͔��d�Tn�E,��Fϭ��ix��E=���/홀]e�*Q���9x�e ���C 9��b�Mp١�QAҪ�'��Rimlc�*�eS�&�4��rh�b��M���/P 4�L9e���B��`$F�Ⱥ�����F�R|����d3T��֨�f$�%F�>[���t�u0�(E�$[R*�SS��R���Z�>����(����ӽ�kB�*s79�f4mF� �9�=���ލ_��ү�U�o�t�~���w+X"�L�K�PZ���a{"g��Ǻk//�9�B��B%��Y��(2����Z4j(�S)V�?IB�<�R<�n�ʓ倭[E*PV�L��c��I@\������i37ܰ���Ub�!��D�=��Q�N�*�5���I��t�.���e$�:��������KD�a+�l�����ۄs��=�۬؜o��j�\<�V�_c��կ�m��v�-���jv��ۼ9��A��鉜-��!�M�es�w�b~�*AU?�u)~��mC`�`d�2YϔVG�I��5�E��V�?T?�u�����������0N����&�&H�P�T�"�K�.�d\xD��� X����[CWag��0Ì5VH��,����O��3�h�pHZ�/�����kQ�Ȁl��a�۴��\p���G������E�bʀ<�>fq9b(4�ƕ�3�9-�^sG�M�y�$WU%a}�R�8Z𩀣<^�6M`�TQ�I�DUV�E�L[��W��J;�}���p� �����Q@�;F)Q��ϰ��0���DS�=�+mu^��ۤR�V���5���-d�	��TL����덪\VRj�s7ડ��f�uw/�=zmj�DX��֒6ڥ�i͙���Uk㜾nt.`+x���-���T	��5 ��<���0���+����p��
z�g�UG6\�%��= ��s陡>Y�`� þ�؆MWq�W�I}|��a��7gW�'�;�P� ct�N���b�w���۷ym�d���*er�_���.��)�H���;����Qxî�xx���"�ݫ'�����o{ξ^�ܲ[5#��Z�?>cm ֭Ԑt����[��҃_2u2���@4�gە����#%�����.
��$�R�Դ��ˀ���Q'f���w�fY#B*kQ�`���[e�b���U��\����dS�p�5$0�4X��l�GuK�+�5��^�~j���U����4;Q�-eW��X�0���+`*����rPM,=.
} ���n��OTX*  I����4?��H�*
e]aWh.V,/z8�&��3,�y�b;ㄡvZ�ZJ�z� g����*K��Þ�h�����.Y�q��ܪ�.V�������e&��	"B`]�`*ew����+���-���{��y��G�n6�Xw�R�֏������m���u6��\+����d⊔ܼ��$����7 ����"#H��B����xEF�v<���t���M� �6E�oD�iE�@����r��5���8V�^�S��6̚�U��!$�D��T�I�H:�D�A5O �s*~��<ʩ�7�H�#ADXk�ߪ7���z�a�J|׈Z ���Tg7^u��������Xo��r��Z�k�\r�5��-\Qg���8۬�%�DU��;^!Q)��-�&1A2�]́v��>[�i]~K�4 �E��c`�/�}BH�ܴYD��
4��1c[O⪹��p��K�#A�WZ�?���_�$�R�@�%���v�g�ұU�T/�����ܝf�2��ц�$�e��{���(�0ΜT�Ï� +.�x /e��̓2���K����r0ab��)�w��1��{t��
m$�Y�cq>#O�,A��B���w��p�R�J�5��9���Y'�����h��{��aG�>{w�)�ϱ��~�N1����۞��l,�$d�$`�{�8���UW^f��K��'�
�q�a)�"`ז0���ο�"kF�W~t�0�����X���{����6��<|�p���������W^m��y)VE�{X���m�?��hP��z^���=*�n�1���H�ϟ[�Q�M2��s�Av���y$�N�-����9����4��O��-�ˋ�얗��X�����F�_�i߾����]�T���� �9�ʠ��0���L�0��*��<��K*_60m���*����>̎�KU��c�(�z�y�I��no�G��m��e���,ꔄlY��U0�lվ�6�^j帒��@���k�(dT�<!�>��^WS1�,_��8hx�RL���f�nS�z��%�f����]�����6��3}���*��T�W6��8'���¤4ok���ݦT}v�_�3�2��Cw��jD��������X�;�\���b+p/��n���![8\a�&�B����%K�6�@>�
)g��k�UJ��1�r^2AN���NjD�L����qP�+���#�Ęt@�U�F��x��-+��~������kKԪ��X�]�r��z͌�9�����~��{]��Kϱ��^�D��#v�cl�IG�˓��CO��ڋ��ԇ�>�&Ki%J B�*VpMY>f�M�<�m�*o�>����ۄk%VIZ�X5�*w�=������F����A5L}-°�
X��z0��rl<7���e3צ- �"���ʰ�l誈i��f��r�
���#Cl2��E=~a9S bj�IC�t�W/(�F�2�щ��H�5��9��"��zU,�e;�c�V�?��`���ǖm�f)�������#e�X��f*֙��� �
�;+�Z
�+��'Ӫ�zg/�GH�
\�rm�H�F=���ժ�`^?��*��) �J@�
�d�bO��
��#����Un��El^I!��;ɦ���4ʹ�W�VU�`�x�D<ju�Xz�:�R��ڒ���=�$�5ǁ�ށU�˺�����5����XOu�|�������(D����b��y�i���]ƴ�_[���zf;--`=њt����r�x)XE�*i�M��bH<%e�r5J<uED@����a.A��+2AI��h�,�O�~���u������_&����O�9��=�>��g���=�@m,��'���'�.�g���*:t�=��|��?X%!��k��N��s/�+c����m������'���mr���XÌu��7�ԏ��^��S�AU�E�n�oJ��ڶ7'2Ttٔ�#ޞ�p3����6�L�3�H�3\�y��#��`J����}�
]���w�1m9��u>!���l��]��TwqxħR������)�vХ�}�5%8�#��Q��2ѐ��h��^�}���%h��WB�38F{%����/����/��[�[C�Q-}��JBv�&���U��uU���hb#zg�8���^C�����B�h���J>Q=w��E�U<�D�Q|E�M�+�_�#XD�r��eJ$�q�΢9>�F��Ɖ!�{�����Y��|2�k�����Z��7�X`���I�ޒ�\i�T5i�߮��������U^�6c�@�a��#�,�	��.b�+0"He��[S��x����X�:�k�3�6�c���[�>pr���2�R5I��ZEF��ȏv���q�L��^�M��d���/�\g��B`�'�WU��2�,���ST/�U�ڲX��D��c����s����x�#�Km�'����u�3��������h������Zz�$�W�q���^ak6;+8��0c�>���5��sv�y)8Z[:,6��ж��=����m����j8��@V	�� p��	2��T�2�綽Ԁ�uϯ�\�u�g�JfT	�Q��^T�����F���B���/���D�Ȯ$�D޽�{���ny�6x�>Ϩ�$��
3���*ڰ(�Z?>��;)o���26ͱv@F�7?��� >F�m��|3������܍�֡m���H'گ��c���M8�^��z��Zà@�Y��G�����,e	e�f�YaQ��z�]� X}�ISQ�����XՆ�W�1��{fL���F+���PzV��|��7C.aU">��XK�C�[��J*��I���Q�Ҭ�Fs��pSz���J��� �2�̇jbܸq�����(!z�($3�$4���b�}�B�m0������a�Z�X�8�X�+��ȶ��ۈT`FS�H�Yx:���B�M�Oi�>O�P���U�T`�0����$iF�����\�h�ai�L�#y�rVay*x`ba���@�{�v�  _�\��q��h�Fp�`/�K�`��s�mm��f�2���}1 �/`�f�e�K�[=V��X�=���J��X����Rp�ZP0&`{����X���wI��A�p`�XT� Xӵ-`&e���� ��>�O�O�jS%�H�-Sp�N��}$--5�����b��%�û�WHl���C╎ɥ���7�o*.�
M��~�ꋅ<��a�����q�hVpui��h�l�]t��Ev�k�R�Z���h��JB)Gv���񶦠�~u��?�x��8�`�;i��ާk�L5��~�uc��ӓtL��i��m�}�66v�h�b�{��HD�'u�?�t|%w���<߾z���[��g#��⋬C������7 4�����-ߗC$(�t�����N�f��E�
�����^�)J�}����|��*�s	D8��NK��^y�;y�1�v&i�m�*��}���e�~�a��۪7��
p��#,w�,`m��ڢV	���k��~��(7�s�=���~���a$RRN2�*3���_��V�.�~�~v�I�]��CL@�s�%aA���ڈ�P
.]]o.�J(M��SHRe���	�8l�h��VM++ͯ�0���2�X-,��RI<'�4Y������Qĥ�A��*R7$X�(<��*٧H�u{�9��)�������mK�_~��V�=��Xu�[��L0�3��
��U/�{:�/��( �*�K����$dS���|����u�VdHY��B��͸�8�Wbms�X/nIMq ���R�=�D��NpL;�`�_`�{���ʬ5*X�q�X��)��S�mTz���wk�m\���+r�]���_d=[S���&��p��7�dZD���2�clua�]��'l9n���kD22:��E��^�k��AY��L��*��U߸�2<����ؿ[���x�Rr��^�N�U�� ��6���<w��9g�e{��i˗.������������T��c�.��f>92�h��3[���윍�H)XzV/������Q#?�u��y�*�t_PQ`}r�U��m�v֒�N/��;�"��W�`l�ˉ�`~�s���/����6g�|��[��z�����NA��'?��>�̺vf4�s�Qe���\C�q��r��dk*OUV��|��Q�L�f����������	�X��R���}��O�u�y���j�T�+��8��{��(+|���;S��zzÊt$m��
���f{`M���q!�plX�Y�sg�qV�z�a)xww��M-�*c=�c�X?��'{�u��ڮ��p|"$/������� E�,4�?��o��ġ��T�R�ޥ�*�����Ӂ}���\�Y�׮�q	NH�B3➭F�t{eD��"=U ���۾v$�'��=����� �y󖖝�m�Tߖ/_n+W�ìYӐ���j�;J��h�s� F�Xs��ڭ7_�)�ϼ�,8{�F!�劘S�ڕ�r��|�U0fsí���\L*�?#�ĎVY(e�wFg�����
�����FT�a�b���m�l2�\J&�I~���ƁU��AH����$09���g�b�RkD�{��Xw<�a�����#�W495XP����k�~����z�,/.jf�?�T�"E ��+cU@Z�W=���X+���1�mw�9Ζq�ƽ��t�y�v衇�2�i&<����wk7=RT�(�`Kh�s���[�nem:��C�X���kc�ŹI��VH6YÅo�,�~{���gx��o)2G�A�I7^{)e�t����J_��N>�`�ؾ���5�q6�A�`��<9�	ZdaAΟ��^yc����O�<.#y4��5,g��|}�Qv�I�y�t�p���{����3�X\j�ա�Q�M�C�!�㫽���Us��M������ofۇS>U��{㏿(��/����ԡC;��c�ߊ|?���`�?� ��jx�%�d��B�ƨ�k�H.�В�6��g�\m�"4��(���9�e���̙=��o��&2�	��2_M��T9TW@L�rp[͟z�X��Nb�Y�ۖy.|ߥ���frCnA{�2�+�T_%=3�c��b�]�w�l��l�$��\=�R�m*��q[,c��{��s��HŶ��s�OOH��[�Be���R��YR]��}ډT�R����av��j�Ή��V]���֋у��^u�ֵ�|*{��u�����~s�}��R{��g �1���N%����9N�1ƒ���:���t�B��31k9Ǻt��u�oO=���GEp'ğme��s�ܭ;dڦ��6یY��ZI�m��FZ2nY�X�ق��	/��R�� k�6�o���+o{'��~�<�$� 3�Ǉ%�"�O=y�{�Y��9���Q#����Zm�'L����h]QE�\D�"RIwG��"q�9\�Vm�z9e%�I�
Yr��SK��M9�Lty"̋�>��ki��͝^���I7���~>ʞ|�{������eݻv�������IÆإ�f_�)c����Z4϶3N9��oO���r��ޔ��G%�O�#[�¼�v�~}숟�g��Xk�G�v�W�6��v#�udȕ�6��������p�����-&�}J�z�j(%�"`q��[!T���Rp�3���ʏ5�p�m\6+'� �H<Ěf6u۸�y��`�B���b�q߽�5�r�e�Mf&V]CVPj��%6��|	򑖞�qr�	m������dh�r�	r�uM�mo���(V��;�J���1}���<���<|5����-����[�`������,^���/\�4@E�ޕD��LU����+5��Ū�7g{��Je��|_�`�v��3k�I	���qJ��*�9t�>��������[���v��ɓ!�0��(�=��	����z��Ƀ��5������Z�=��c�7qk4�k�{5.貋��$hOV�Cɶ�L4)9�� �3U�Tx.}���L~���NX���Z�tj)�/!I(�n�զ�yMFL$9�#aI�z���ֽgJ�X��d��ɧަ��xIA���K�R���6}��V��ā�쟝a}z�e��ͱ�{���b��4�Ð(�=���6c��	�|hM��X�
��#,u���J+h�R�2֪� �� kY-����+7B�"p`����M6�}�K�͆e[o���S;p����!*�������~"�,Ϭ�- ��ȴS��ֆf��ƱA����~�XS���Mu 3�E������+.8�>~�s{r�S�|�%�]N��n��nˣ?PG���X���� ��,��;�����EJ
M:�h(�`A)�KW�z��V���.]��Q:"��FIH�m2���>��{��͜��^e��g�̙s�����z�z�)R��|�"��3    IDAT�+�l�8�d���'�O�s}s�BA�����۷e<\-��;�b��ԧ��y�<ـ�i��i
̤���k�1p�FpΛ�!�� ��x�~��[�������.9�}z��R���H��Yff�"���m�)Vp�f�Z1�Q ��ܭˬl��`e��##�S0 �ѳ��Ű����ZUw~Č�s$څ�H??;
��;�;-S3��c�6��j�?��p��ΫcW���eRj�0�A�w��i\sfͱ\�T��D`B�����s��$��(�5@ �@,��!���.�$�k�$a��w�$�T�iC�B��|�ߺ0�)�eR�;n�g~sU�|�@hbo�<�3�X[��]�7�~�8!=��e2v��<�|�)���L��T@�PKKӵѾ�X��> �����T��;��U�7����K�]�z�]=T9�w{�n��{������}Ħ�;�n��I{U��ʪ ��IRw��R`�@]������-6漢�~�R����/���k/��y�׶ɉ�)厔@,�4V)ƌo}D�e�mI�j�WA�A6��s�\Wǂ��duل��}(Rj�,"v��^��76�C�ڮ�(��\��(%�#c}[�\�]t�Ev�1GJ���n��g�U ���t����/	��]�{��z c@���뷺�vp���a:�JF��Y"T@NVE�n��6Bު����h�}�׾y�=��l����א1����ѧγ*�|�p�Ə�d�~����[eo����JaK��Eh���`�+�g�B>�����؛Պ*�$��1I ?�v�Gβ㦍�&����/���[�Ѯ��2;G��G�}�n��!�V�rY�� +�־*IÊ[��[!'���k^�rV	,�� U�zQ�ӵ���z����B��Uw~D�jΑ�e�"uzbܘ��!�<.�\��ޜ~c�Dk!JV恌�����e�a���2�z�:8~����[o��%˭g�d�HԹz���E����R�������di�/���)Q�Z�"O1�@ ߃p�Ӹa�ԩS�{���@nTNfKr'�J ��[o׾G���R�^_' nk��'�����L�Y�6A�x*�٤C$���ku!����3� �p�țd�d�;*uwe8`g������N>P^�������H���B�E)V�?j�L��Q��Bi�"��cU�Z�~��>����������n	�̔�+$�Օ�Ҍ�b=z���U��%��S�k��s�{	�	�/P��s�L��kl�s���o���n��b����Q�Z{�w�X���UZ���C�>H.>� d���������� DfkVKy�q��'��Q+r�m� o�Xa�q�f��p�av�'ϵ{�~��b�~�8������ɝ7]ҁ�e��K?f#Ub��n��ʞ/���G?|���'�_k��w�u�]�W+�̳���6_HNQ�)�%��`	�C�z>ѕ��v�i'��h��y�#�K&[�z�UVU�؉��o�<6�~��GU�{Xc?��Vz�g��z�6m������
n��z�XS��~/�f��d��A�Kz��q�X�{)8uT�xYYY�&575j���U��\4d��'R�"R�F��S�`�{V$����r�s��q6w�\Wn��
P��ă�T�0���=^ ^��=�c@��^j�/���p���&�ۀO����>�'P��K���n��&�&���`�=嘣�ȴ|��0���Qּ3`u��X�X�].iti�aPi��x���KY={����2J����2��=^�SE�}�{���r#���Z����v�q&72��E�<�3jc�.i l*�bE*�V�`����<l3�NX��K&ɣ,�q��O�����<���>m�+]��{�W�{�چc�v��u��=�2�'Xﾽ<c}g�R��QKi�)��`���ҏi�Lߏt��<�)#��~��V�+�J����u۷-[����x�و4������rR���/]����{I�(?�¡�!#_ �\-�4E'������7��A��k��y��~+�7X�ЙV��¾������}�����V��q��?q� ���@�?+e���?�q�d���^��ҋ+j����A��.⒋J���3%ix�1�&Ms�23��o}���?a=DSfCf�7��Ub^�f�D�U���C��H,���*���_f��V�H#9]��kn�W�򛒌���W��"+Pd�D�����#q��$��������W�Ք� V�Xq���5��(��6���M���pf��X���T@����k�o��1����>��L��1�[�=4H��EHѽ��	 ��@��� ��#�e�P
�����S�w��1<��� W�5�9�(�L�۴mv�!�X��P��)�k�X~��e�>���a����E�S�#$�U�U ��;��_t�����8G	
�lʣk	8N�����K��%rG�*��˕��>j�%�T�,9]ә$,�Č�y�}W`-R��O~�S�u��K��z���;�p� ��,��1t5b�*���W���t^���v�.|��5S��I^ ٜ������okݲ��͵ڧ?u�9�pP]P�������*��YT~>DyAȘf,������O?m�W��Vp/��}�
�l5�j����~����W�'k�{�m��<(�r	"�d�̰�j�]�ѳl@������m�3O�l'L�j�?���\�F%�͵}��KDo�{��ϑ�y,���� 9A!�5�5�-=��T������̙k5����(�ͶC�d����7�f�k͘��͓0vvDuS#cy�R�M_�N��~~��1Ie�t/=���N^����
N VXk��%P�ܪl,[&����:�n6m����êk���*z�ƈmk~��V���� �v�ձ{`Š`E�F��a#�<�����1���'y=J�v�ټkU#��jI婔�{�E:�-��r@]]�%2%�	q;�һ�:kY�0-�i�)���쬭 ���D���O�2�V�X�~�.���svQ
N��R�� 6e��Kr����(Ȑ�H��n\��8I�I@�&���"iJq���}�-ZWfy*M�
T� ~v0�w�[��h&Gb���BLdԅ�06�S�	)�j�kB�)(�%�J�R�����-��=�m���%v��q��x[U�_8s��uǥ�����c_5b�ׅ��k��K�9��챒�����F�B��Ȩ��' �X�y�ꗽ���Ə�K]�"�|��. �Rf҇w�#<I�U�D�3u�5���m�03��eG�y���R��(׀o�@2釨��BJ�z U��)��K�9]Ҁ�[�lX��i��Tѷ��1�(�z��(�4�:ގS"�z������C�D���+\(Zy��Gu�"�6{�UZ����Vm� N
!�3����TD��Sx�/O�:�U
V��I�u��_+X����۲K�P�w�\W2V�/����w� мw��ݺ�^oDn "[DH�r��s���c�6�B�8�x+4J �^�z4���-�w�ή3V�a2F2V�ކ��J��*ec�l��7W���N,�4i�+���j����T�e�fHKd��bPA���q�J�0�yi��|n�I`�=�I���KW��U�%x�Jd������2:�c��A.:���V�26�Q֘���L�a��:����h�ڶi�2a�]w�?h&���u�-]��r{k����kY�r�O��PF��9G���P I��t�;�U��X3��'���Q�+?w��1R*��ꕵ���i�.���p-��ֳ��+Wi�V��=���iy���x��{�Z��X郆}�X�ܶ:{M��&e��K�3/K=/;]d�) ��������׼+ڼ9 ��AT����M<�,�j��j���U&e<E$Օѻ�>[��3�� YV)��i�H3ǽ���*E�F��stḑZ��͕�sk]�~/�>�N`��C���Շ���Zݘ����w�/ZT��;�o-�ϱ�8%�~�^��Q?��=��Q���쒋γm����OYV���Ti����l[ّ�B^�ּ��ets1�F�5MTB��"��^Gw~�Rp��M3}}����,��)�f��� /u�ձ����uj�6Tuble��	6c��@���E)P�� "�M�"�H�-�Y�9v�L�G�Qi�БV��B�Le��M8��ˤM�Oї���ιY�n�<��=�܋Rv���a�qN���N�4I}�2U�TKcv����n�$-�4��4���5U��S�ԪўLe�$�-誋�T]f��n_��%� ����wۺ͕���@��+�;֎�SR
��1��ŧY	��3�X���9
��z`G`u"-a��'���+�U���"�2T[e�<��K���uƊ#��nش�^}�e��k���R��`�X������=V���&o ��+��,�Gf���5/yS�-pFi(��8#���;��)>���I�qcO<���<���ԯ��RKl��G�3���'��q6�p�<�w�K�=V�;3q�!bݾT�����v�>�M��k0τˎh�{Ik�.�m\{���,�V@�ۗ!c���@*M0!/�����UoX�H��N�~�"�:�V[�b��>g��aec*�S
��=����� �{��FS�����G��&���k���?�d-w�o�gs�c���cmn�0��O�X�ŔQ}�j*7�`�������MR֖kE�fRv9���O�v^��Փث�Ay�m:�[�~ƞx���w��I5�V��y�6y�d[!>��ի;��IS��P;��Es��B#���
�5�+�
�mJ>j|dH2V-��fl�tOI��w�;�̓|.�/��!��j����>~�%kO��⾅�=��@r뙺��v�g���36~�G��m���\9:���-� !/e)9��i6U>)m�����]���cM�M2/�qw�F�֯_k/�:Áuoz�����}��7����f�%���\��Omh̐�R V26w�S&���6�>�l��s�z�J��Zb;Q�7�Y8�Ｇ��-� P(�v�!GZɠV/�kV�� �2�A$?>�@r�-����I/��3�O��0鱗6��Q-<'�[ �x�a��o�`q�宪������K����p�� %��&��fxE���Ys3��;�k��TR�Cx�`.���2�Y�d� kw�XS�Z��hN;�4�1�y�O�8�J���X)�����`�U������	Xkk���m[4�1�.��;�����#���Pն&�V��e����ѩ�%�D�Ԏ/�{�	�D�5 ��¬yo�;��H�N@(R�*v�
V�5�{ǒ�iS��ƌ�q2VX�� �4�?�w�}��OZ�ذ3$	�j�[��̪Z��+�J�HRM�ؚ"p��/�L�|x����-aP�sd�p�$f jj�{�	^�H����:)kV�K( ���Kk��H�*�^�Tmُ�c�W�=+��q��b+�5�p��{����iy������_�o	D �y^���H�{�$�b��hr�M���g���������e���>�E9�N�8Sj(�"�(f����x��2h���X��J�.�xS/�g�b�Y�Y�P�-p�d u�#'摑���ʫ%�
	������m�R�5]d%���؅/h�"�8>�\��]�W~�zJ�0Meg���/��`���P[UB�Ώ�-��Ⱥ1�w���8�W\Ұ--�K�X�c�
���<��;u�{Q���ݱ��"_��z	�Py���^i��Qg[��Ξ}�/6w�"+���H]�!�n�ZN>M�=�@�L��d;�X��3�1l�|f�݁uͪ����h�̱�,cX#+8����YWa#z�?]�=�J�f�U�r����\l5o���Z~I�%�p�t~I��� p�]����,:��*%s�#�`mR��Ϣ��{媂�H���RW`��Αks�jE?�<YH�V�d��қ�1y)�4K�g��4�C+ɣT2Z�uV{�
�nz���t�.���F�k`m����M
y�T�w����#��_�� ю~m�|Yzv�х�·��%ԧ�Aq�m�E��bf؆���>�w�@�p`Ά�� �-Xc�v'b��]����o2֐䒭������T�f5���݆�p���F캮;�X/���
+xѢE�*F�GW
��.d��kVgL�&�5�5�O?���������4�'c�Q~�|yS����S����0	�f���;�E+$�'2K�TϨ�5��bI�~/���{�K�����f�?m&�P効�4ei1����&Rю��=�ߗ�����
fU�s�6���iR�����2/r� ��ח=47�Y��e�h�
[�r���I	��fp�xxU3��$*��:HH��z{���������D9g�Q���}ܦ�i�t
����Y�\�4)/�|�^k߶�+�%���V2_��)��	R鎁5��z9�l�=y�UK�r��m�Xyǵ}]�K�y���u�� �� ���X�]��Y�w�<>�8���g��g�E��^�H8zI0��ŧH��6�� =�\c?6X:-�8ܝ�wy����j���	p�H;���鹆	���@J�Xu�P!!�5� +�g�|�����z������FI�P�������$7##g�q�G�܌/��+���Ǌ@�`�5��N���'��;��)SjƀCc'�3���|֎��C��d~�G����]��`�f,�U=kԞ�f����6e7���߁ ĞD �Dd�q� �@I�+<i��=���M9�g��bD�3V��� k��!��KH��C۲�S��T���O}��:�P�?W<	�O7����Q�S�p]�Yo�����{[�M�+B�<��Xf}�4��ud�z/�nOe��"fsc��N��u.~S�S�7z="j�i2~D5�X�J�@Dֹ��JF�+]h�D	���Y.۸F?�4�3奰n /���V��\K���:��g*c�c�RV�SO��F2VoFn�c����=)I�)m��QBuI�f"3z���iֈL��?���j�K!�7�64�X]��Kf���n_��������/n����D�T�Q�UI9Y=V����)`��p
t�r�}�p�����J�z����Jƚ�'�J��99����Aj�@��M����w����%� i���{k(���[�$z���~�G�ܨ1ce\�k�� �nw�t������%Ŵ����>c�e�͊{����/߻Śs�Z��?Mچ�f�L�%L��5���mg�p{r����#c���A�j�� U�F�W,�(��s�	y)�X�?�������5X�Opa�`	r��K
�}�F����)�����w흷�H�h;��z�C�����ݾ��;l���mvX�����
Y)u���6�TρC�ɿy�J�Gc�6��gِa�T�͓%�������H+[:J≤!k�4D�R��gvw�����*�F�K/�he�7��Z��]e��!�Z�͕���� ������w��{e����j�(!��.r�U�=YG�?�I@h]�5�N8IMgC���Ϣ˃� : <�1�,1ќ����
���	)G��JY�RHք��ec2���2OnVC`�����׈tG�����8�����f�k��z%� �!{��B^�t�c�{ V��;ph�E`=��3��d�{u���c�kj�� yi�o���_��2�Z�~��|�`����^���"<�����;���V�1@�Ax �K�G
�ؐ���슼�dL2R�K���(��)*|$�����k?XW�Z�=�L��<��5+8J�R0�6AО*��p�WC�F˗��?��|��G<ӕ�:h�ƌT-������|C�����5e"{�	�R�<���U���3�S�bz��'b(����SR`�_r�4��͙�О�%���T��m���:��(��g�ρcR[f���+kVƊV��W|�ƍmo�����Gm�ƍ�#ԷNYԝZ��8�j!A�(��Z�ubF/�*�`+`���Xw'�gw�ZV�>ŕ���c�AQZe_�?hb;U�ƽ.y�xai�nﾫ���h�$Ҡn�櫩pP*�����b
�%����@B�DU�u��R���RP��|    IDAT�c��	�)d��E�BPç��K|��߇��s�׆��K�p�~��J����r$V�.c�y	`u�'ku�Gt��;7�`�R
���Y3���J)� y������lG��YU� /i��?�o��!'���aVI���A��/~����ϼ���R<@���V#n�sR�q�\��M��j�b
��:W<�T`����vUbphb֞}0G�K�u/�ꩀ	� �Y�LѸ�T�V��@��;o
B.�ŸM�V�O]@�J����4�w̡c�	��pͫ�M�ƉpN���d�Y�J#3�c�bE#�#�T��T���I��aGP�S@��Z�z�7�<�`�`����g�n9��η(#�7���Fe|Q���$]��S��SP���:k�,��S)�Q�K�������ÏpE����'{$iȹ�(�>��i}����Ų�f��ƞ���֋�����Ӧ�h&PN��0?���p�i�
$1H�8{�]�=-:o��I2�T?�X
����9�y#��]q�g�p;Y��v�����AB�`7NG��w	��K ��?��Z�q�
����n/�ذx�eK�i@�^�)�Ҋ$�X�`f�̙>n�'�&$�2�ا!f�`����~��)���Ex(�k�kK<�m���`o��w��}��
g�z��7�((�j��*�
F<a���m����o^��3���g��o��Nۖ!M��>��)F��bi�gI^U�'!c�B���;��$Dg���,�$�t쪡��2�z���4j�3p�)�|Z5�z��u��X#�N^�+�8^bg�`�|�ϱ�J�`�=H��,������[_�Δ�9�K7�/+wy�wP�R��J,�Z�d��*�cf48�%�,L�+�7{�ѓd�y����pUS�����|%�&͘��=����~�r�i�'�x�ƌ>X8�k5�����m�J����=ҙ&%]>�#�'��j�������y�r�����Ϻm"�w�u���U-|W�2\�©�#f��q��fo�mv��^|�<��>}jS�Ԁt�� �������85�Gnm�;�x�v���>	�)0s�!)	D�������p|�;׌����v>�2��}����&�������кA�$�n\��sk�W�"���íH�nw5��}���p��Qw��#�&��Ȱ�O:�$Ng��O�?k�?��+/��c���g��� ��;���>ޚ��s`M�wd�! �Q�l��پ��١�8Ȼ�_N�}�s��i���Yc��o���\�Y����U�	�}��V�����G@ܚ^���Ӻ�]�}�xR*`@�������ƒ��f���^�ˬ�WE,�R&��c�|���JpHqv��6`�L)���D�V7��>s�ޏ\��[���Ez��~�۪�PJo4��{P�§���:�͏Bfm�5��LJN=�([(��Ç[�ˑm�&ɦ��6�����m�����m�8a�]'��L]�Eo�c��.1��q�-�{|ZB�eOW�9�����ݏ�v�����M�\6�R��+P�;�6���cŏ۸���)�j�*>���z��Ѧ �n���de b
�0;z�!w�Q	do�Ȯ=��Gk��a'��a ��{���w]�eǀ��H��߅,�-��TY:릥sX�3P8ǲ��k<d#y�q��^
�9�Q7q$Ię76�1W��S�,U�ɀqnW����`ݻ{�����k�b���3�Y�X]���T@����Jq��g�b��x��&�}y�J������kɕ�a�zpz�a�g�&͑�VS�T;w��/�:Wj�/���V��Q����[M��A$)�)X�=���Q�>u�X�+�*�ܠc/�6�p}w�6�E�|Oo�'˴:�R�+ϣ@*[$��i٥�<��R{mWI�A�z;�cnaH�� t��*�7JנO���|F>��<�u�z���ԥ���3�<o�ǌ����m7?��۫v�2�����~y��.[�e����	�/��:�����r� �Gn��i��fZg����*�oM�B�{�K�.v~2�=�c%07������5'�O9���}}�����)��ǥߤ7�3��['Xu>og7��X����mr��L5 � �6�*��a���!����~�F��;+8j��7t�!o�s~�&���"k�.�쾣=c�L&q c}������5��4I�ICJ����	�2ά[I�1��mԀ�^�����F�&>l����̟g�\�d�Eۨw��v�I�RR�'��>Xz��?��P��T�
�'O@Ɉ]^�t9b��D�36�ێ;�X�%��>�N�p�����JEu�+�O��:��zO� �zr*	�T5��k�߶JIͦi��{�:n���f����=���ZY_�z�%"�~�Y*�������~k�'�
Ln����^޲?�������i�����=D�z�m��[��F���]j|T��T_f���~ky)��!/Q
�������'�V$���!�ɉg\�=�Ό5]�f�ԯrs_�7/'yeǁ&-^��î���t?�����N�T��3� )�_j_����n�����︷ڕ������z="��X1:G+8_��6���`
�=z���}��|�
���Ώ��B��"�YN�G=F�#���k#�ms� �9��::8�)��p��5��Y|����2'��Ya��P�6��#'��.>�9�3W ����6l�fk6m�u�V!5�*�a��|��ur?���L;V�1� ���h��w�ɞM�i�}��fG)Xf'�N9��mV�^'�+b4 1���K�����ڕ�z
஻��[WGI�U��9w(��p���r�����t�Fe�E�+����n과L9`����dW�$�kTBٵHNA�|5��4]6�g�t����������q#퓟��.�lw�}��dP��t
SZv�\gt�3dt>[=V�X4nC�`š&d���	����n��z����kz�Avș�#`����?���wͱn�*3�q�=���2��$z�e:J��zo��O�*섡���G<)�k㍴w�����X���V�)	?-@z0��3(QctN�5[=!�Gw�������C���%ZL�K4`�נa�n�(��"�������g�.c�7=V�od��X���Kk����e�O(2L�f#�7�N�z��8�(i�E�lC�_�(��NJٹ},��,�p�vvA/�P�y�kU����<nO�<���5v"� w��k�M;�H1�Wz�5#W���[��
����[ns�=V"|���+皱���_���k~t�M{Ӑz�y��
S$S:��Uv�}�c�V	X�1�~'�n�.�R���12p�[��f��\�>�������!�[4g�C"��z�0͝6[�4���a��nt��
�Gb�N� Yӓ�fͯ����T�R�:��4�,`�<v�`���!{��H>��q�d�ñ��co}��q���{�c��~��M��
Xc�3j 1%"�N¸IT�����J5K�!��8��f Ou��Ϗ�����x7�hw��;�����������L�]%�$ ؎YL�z� k����-Kl�*Ѵ�A'�a�{�cE��O߁Zкf��Mw�.6���ۆ:4G��5�DT��s���q��R �� ���
�[��=Vz���������T�ћfU�J�5��X%��M�S��G��GN��}zi��f���<l���R�hvG��Y�������'_�#�� ��s�L���N����ٲd�l'���:ǚ
��5�6�4���_��D*��/Yf��CW��J�45�6��%P-��>��?C��U�^ �tEE�J���~<�� ��m�A���� 7Hn0[�f<�[��x��N#��vA����<�۶H��A摩"�}�	��%����M����+�]~�+=�_�{�Q��w��z-A�y׌�Q�K{S
�`͚Ҭ�$�g�e���i��W�N2��9��.�Y{z#����F,�)S5�Y5��*p��U=�2�2Z�;���V�6�l�p��Kɭ���S$����8+����<El�5�>nSTT�`��X�4�{!/���q�شi��̹���dX�l�[�bܦp�H�?����x X��|�=ow�����@��گ_�0n3wnG��A�&�X[�Qes/�O���u"����/v~���VR�g�E��<�E�;��2Cp��wCk�w�Eh?���k��Z4��3l���3
*��P6���`Φ&����Ѓ�:ʘϞ��!/E?V�i`3ns�U��3�k߼ŝu2�
�EtґkDw��q2�چ�뺷Z�Ȕ���n��A��XҲQ��]�U�%�սJ杩�&J��*��,�R�z����&�I�2�H�h�D��	s|�SR�|��PR���=��5R
N!/1�z�}��ޮj�F簡Y�e%2o��Ÿ�&�,K����ۿR0�q_��'751�����=���ji4��2�]�JPi���} 8W��E�=PTP�|��}����F�5ݬ���x` p�QS-��`�k�"U�k벫kK��ݰ)������g�`�%�UЫ`�%%D��-�`�%�����������鈎�����y-ʘ�0YxDJ��th
T$���V�y��%��������a냆�rq�&]�`x�?����>7($J��#K��r$c��R��� �i|���[���m�����:�F �&���k��w� ٻ2�'�S�ݜ�h
�bl� �Ln��]���*�kR����Ch�%�I@(�&�3�ԏ2Te\%�D�i�aC�F���2v��e��K�5Ǻr�:��=�dof�nQ-���ʾ!��uר�Ym���nq�J%���E�H�o��֔�ā���k���t��?l�翥y�R��li���u|��3�_eaY����������A�'��u��w�:�1q�}xn@����cH�*3g�F����^��x!�����9���S�KEť���_n���&e�����M��j�J{��.iج��=��^�'�4�OiIq�'�/2�<e��_x�V���`t�>����fN޸�K���;�0����"���P��p�V4h�\D=ןxT��b��n|
Q�J�'w� Pn�և���	م���y��#)�XY(�0Z�ەf�~����ZmҠ7��%ȗq3�(��.�*%���־m���ɐ��P?v2Vf�Z�b�������{�1h�;�=�5ĥ�Q[W�j4�-�P��x�!a��t���������V��i���tVz� k�3��*C#�M��.$�&w�g1WR`HK�I��wV�����%��U����Lv�? �]{c��5S[�5�-%�&=���z��Db��3M�6��ͮԸ�i$�gJ���¢��λI�T�s?��J;H^y�}�����w�K$ث���B��y�pB���U�r�KWA `�q�>s*����ީsB�����H�ÓME8���SH�9����^���$"�'�,}ue�"���Ue��_��&�8�V�a�q�o�~�c�RB�%��!. ��j��������-r%�۸������O�7��Ve����:u�@�����k����W���-�!��Zv�����	A��{�����=�#����g��!՜�6����9�*���.����(��8@�{��TР,��") �d/��P-aySf������ )� ���r		����k)ȏ�a�;\QYn�����*%񕡛'+䥬�Ş�2�
��k�w�s�Ko���͜5W�<^1Af��{g����GD�aذa6u�T��$0y��?�� VD��c�̸́9��X��?���R0%�A�9�ΐ��W<$�GX�H[n5�� Ì'���>k�B�l[ B�!E�$@��J .�EQ8�a�N���})`NT������!R�ֱ䩺����;YZ�(/	\M�Wo�L�wb���݆���D�*_�K��U�\.��W�G��<Z���q9��ww�Hzw���))v���rM��]�DH��`�9=`��\#Ys�^	@W�A5h'`%Ӧ-(`ո�����~�2?����^%R`�,!��,�h��
X�(�9¼<}��d��Tm��-��쩻� k��U��d�������.`�����լX�h�����Pt�7rM&�#����9Z�Dd����O��c]`�Za;��3j��h�R98C3N*�4��j��憲M������وL)ݴ���%0�����{���̄�Ҍ�D����Ǎd�����O�'(�m���]x�U�o�����e��y@^*����T��M�l�Y���
��Ksu��Q^z�ŗ] "+�Uˌ�>6���|���,
y��ư�;����#����L���<�!�oLǸ�I���O�����X��� Vzx�dT��HK�尩�`#w "��f!13Ï��U_����oB8܋A!.<���q�d�"�6=A����(�H��T��dI������|�^e��L�R
�Z�(ㅤrW��?� ÎD�3"�!��8iY��%�n�{��C�|W��L��x/Z����S���ˑ
�<%��C�G��zٽ�;�\D	��)x���t���jz)���g��^k+�V�9,�Q-��<���H}t~<��h��D�Mڗ�E�����ﱒ��5�Om�ԋ&K##�E��9*�X_�1�]1�r��v��^RY�d�7��p���aa������U� A�\	���&���ukl��-��aG�a�=p�mU��U�:�6Y��g鵈��h�^ hvs�)��P�*��� -eC>ܰP�	����Ô�)���ϣ��I^HZ|4�[$��,EAn��t���i�f��ͷX�t��)k��Xs�.�-����{�,��}����~�������Ѳ��u��՝�'��L)�r�9��K�l_y�/��
+�kѐ���T�y7X�z��yup`�w���%x�X�	s��{|�W�K�r��Hj�P��);�$�}������������:�U��y�9XS/Mk�N�.{>� J� ����/�no/[�}�T	�P��
n�%~�J[�Vs�b��,��.�X	F���J�򒷡p���}Ņ�I���$�~O��l�[ۥ��Ij���`HyR=؄蚢��%�Dc.I41	1�G"��� �s�g���&��D�֪k����N`;���O������^/(�!�� b�nX���6.x��?�U(\Qov��ϊ\,K�{B^���������-_%�ן��J�,7��.��r'�&B lM�g*�"��Cuu}y�>��Y��@�FV��`�fM ���R��Ҡ��V�xu­*��� 7�µi�R��&���Ubͪ,�����5� �����8 ��[��"��a���]+�EVZT9u��Q��k��J�e�	��24<��fV���Ik�LX��`%cX��/����u�Rp�X���<�:�c�AI�k��o��g������X�8 �,����R1��X�V�3U�'��5�������~��?i�C�QTu�0ǚ�s�l�&�m��������Ѧ�Fo��~o����c�e�O,�]���[���F�H ���m�V0+"����1
�����s�ο��� �B�<2V�RQ���&���y �Y�w�X����E	.bA�6U��U����-��܅r0�Q	��J��Nc�[R/�j_�*�7�%"f��>k�X��6:K>�zl㊋h	r�w]
��b�`�����UV�R�{�cE �te�:2�p7yC�[J���͵6���Y�򹖗�b��Q	/��١���C9�dDA<��Xs���~��W�^���.��e^�mG�:��{����J�\e��r!5�᩹��/@�����-L�J<d�D:X�0���3����>˖�����Q�A@ס��JA"��F���k�l�f����4��M7=VD�˖ϳ���֯O��+�W�>�m�R�_^~�y`�s��m�b���4�!���O>���u�X)���"�D�h7a1����A�$K����|�n�?���׹{�Qy	IC��t̾!O*p�h��?z��s�x��哔Eċ�GU�,�q�e    IDATLk���3V0#A��"��������穕�֩�}����u�r��O�~̞m��E^�TEV�b��@�4��8��{ iH����ў��=�}��RƑ"�2�����LE�iCx2p[�^���>`M�&{`�x#��r�AA�3k6�L7��]��cw����(��l
�:+��M�*�8"Z*�Y�4�!/����^|�y���i�l�,ͮ~� (Рǚ��"�b8*���(��~���c���^�g�ʒ �Y��֚V̕�T�]p�yv�������[nq �d�#R�S�l�� [J3��z�ȳb�"ۼ��Ҋ��Q��g���[��2H`ج�bMs�)�cǩ�0{�\{��?��|dl�u��uq�N�C�8ԫ�?V�X)���Qef��ӝ�������A2�xps��VB�%���uC5��[j��_��mٲ�~r�-��!h��UtoJ�Eի;��ߞv��s`%c�7o��dv�RR��Z�1�T��a��?����6�W=�*�d�4� y)������̡6�s������}�p߅�K�����$�?0hc�%�dt-�������z��=��z��2�@:�?t�U �4r�N�X
M�6����$��\�,&�)�16n��Fx&�6�7U}��h����?���jkSk�M"����#��Ϛ����c�L&���;aܦF"�W)٨���vG�BJ�"��-�
�Q;��>�K�i�F z@����^2C�~+�m��+V[�d�m��5j���"��0	K��P���N�6d� kl+F�[��x	����� h�d����z):!�^
V��M�r��Q/�'��KU.��^�i�t�a�`�<�<h�[��Q)� ��A���F���6�OllH����(i.�)PJ-Tp�����/��j��Q��j]t��4�o�K�ڵkw{��ρ�yb��u��%6���[���V�DZF8VkC�d�?�JNP;ľ�_���ue�]�CQ`��nYg���x�����϶ER6d�]<�X[��z���_Z��̶��w%e!����og�ݞJx�N���4�h����nREg�U���R���n��˒Pu�2-�Xs��]+I�ɍ���K�r�П/^�؞y�Q��Rp�Mt�G�bu��)���7!7F� +�ۤ
D�ir��}�ƻ�l{`���,-���F�Xg��=f���t�8������eAe�'|v��eT�?�x����k�� .왮_M�*�e�d{Jq��#%��;TJN}$6���"��iKE+yy�"{�噲�[����ju1*FO��H5P6혣U�#c]�d�q2�����:�I%������7X�5�v��KY�C �h���ە� �x�	�l�x�#H38J6rڤ�rk�T��?ϰ�f.����N��y_W�@)�J-�B	G��:Ö�K�c%=��b(,���<ɗ�a�T��d�H�H{��-�^*7�e����9����1V�g�zU� r1��0Q��2��4��i��D���M�V��wM^
Ym�4�6F1����n�X���5�X� tH��� !G���X_��+c��3V����v`�Y���Ȼ<�fI�1h�`��.Z �w�e��#O>�l�2V��2Ԭn��*�����у��o���6筥v��XVi_W�?�Ծ����Y�}+]����*��g�G�������l����E��װMD"f�8��X��ZB"*J�)ꤔ��$`�j�j_r`����]��m��m\�o�-w�sJ��g�8-���W�����<���q܆�o�y�Ї|�1rC)�����r�{��MV�QN^b�� ����j�HCr�q�#f������v֠K��&������������w��=�s�N4�K�s���&Y�"�a2N?l�0;��)6|h���g���eK��=����|^���,Y�1K�,0�^����:��)*�\��N�6E��b�Bu��`����{��B;ڛ����{�?lg�:�J���˚m��y˶U
�+T&o�BG�D��h����C1�Rq�n~�1{e�"e��M*q�W�����Ԫ��s��p�"��R���<I��Wl��kߺn�=��?�̹o�l�Nܲ�}��iE� Ȯ������3��\�:}�.f?���u_���f��c��M�6��k�h�Y��M�<�����䥇7ߘ�����^�l��3-����1m��J����E{���v���7�x��;�����kk�Z,�a_��"��-��3/�نa[�7�A}��{߽��|�%{��Yn�<2j�.ל�d��!�++ކ�6V0�6��t���Z�*��c��$N��X� �n�����ݩrL�>�X_���B^��&��H�c=�c�Ƌb��/�ʈFF�*�O����:��`q;�~�ȏ�U�M
��HbۈZR6{���U������}턣��)GjC�?��H��������2{��6�EV&Q���bo!apޮ/J���P-����V�q̔)�:�*qw�ć߹�]��
���~��vX�%���ȣt��t�z݅~`O>5��V��j�z�Vi�Lҁ4R���e�F�i�O�iS��#/������"�,g4�8�C�jRk�U�k�CM*��/�j3
�<4+���I�M��Mלcw��=!��Bys���Σ��`e��I��L���'}W�rV��X���~���X��E�`2VD��&2V���5+�k|t�ԟG`�'#o4$�y�-�\&m�لcO�ұ��6]�6�N��}����������͟�@%������'�{����sz�t;�#�ӟ8�n��w�ڜ�t�,�>�����~�s��_���=l%|�9SB8��G�� �(/�c�)_����aiq�@�<�XV��[o/�y`J���۽K���ܵ�@8����#�����/�k/�D�!�.e����:�ֈU�@�V������1��l��?C ��T4Kk�[O� 1���z�o|Lm�K�5�Q�q�	#���NR�?��k�/IOUQt��yo��%�2w�
YΉ�Y�C-�"e�5^zv�/u���@5�@i5V���<U*c�4���B��ە�v k��N��Z���~�3�I�TF�g�۪l��1�AqU�{�y��}��kT�~ms�\j�ʀ��_�(NH�\��u�g�y��踟z�e�(4J�(Av�8N?����P_V^�*��Uv]���I�g�u�����/��2q�\mF�M7|Tջ{��徏W������"Vn�,1[b���H+�f����X�F�{������'�m+=�},c��>�k_��'7���&��M)85c�])���:b�N����V.[j��� /j���!+=�6l�h����o��z�v��b���-��/\��"�¯��Om��Mv�GO��/<�~��_����z��T���F�+�ڞ��'�ˎ���8G��"M�.M`�*�-R��Vp����>ꤛ�R0*R9*����������������,�Ο�S�ߌr���*uW5�+��w������>�}�F$��*`��=���
��%���d1i�|y{S�e+.�V��#&�񓏲#����
��n�:ꚲz��y�ڼ��ū��f[~�8�f	R ��RYb]3
0QFu_z�V�>���=�)X�]a*�m"�&�u�Ӂ�J䥫�}r�wz���?w%*�r�Uj���h�_ �}��G���2��T��Z�-6�$!j�m�`~��~�� �`�"P�������m�k�����aO����e�7����o~�f���|��y�?��Ȩ�k�Re�>4q�i@�~r��t͖Y��u��XU���5X�X�<�+kXSD���R
��%���{8M[�0�AC���r�
��T�:�&�z�eHL�\�x�I�����.r�U���ZQWaf���0�~z�����w�!v�՗گ��=�ȣ���m��GN�n����'�Wg����q���FJ(M`�ԍ���5��?kvk������kW����{��8�K�`tw�s�I (�=U��S�X��C��]�̱F�`�m�p��6��%����W`mjg>iP���t�i��$�EE	�e�-�2��i��>v�fJ'T����P]E uɪj�3�����͚tP�����Ӊ�d5/0���X��O�w�4�=u�T��+Xc�N.E�3VX�{:��K�^�A�~�3+��?��%ԃ|c��C��bk ��(PWl��\���{�l+0k�RSEJ�ZDaޢL6����TA��Z.Ғ��5;t�@������߾���l��6�܏ء����3���a���^�v�/5jX�B���J��������~�͜���~��8*N^��>%!:�]��:���������e�^x����� /����JI2/�١�<ݠ!�}�-[�BF���ŃX���+̷�i6���ھ��Lb"e+z,ʩ�/��nʵ��G�����4�Ҧ����r��߰�i�X"��6�o�C�Xb�lПlS��WV�_X�XY<DD`E+8W:�(�pCa���RϞ=Xa"&Z��=c��
1��7n����!��UmC���K:�
���y7���X����G'�/��2xmj�����K
�ە��M��Q�VM	<Q��?`�&��G�ʠ ��&��e������L�_��@�T�z�mQ��A]I�a��L��22W4���t�e�Z�(�S�c�pb�6����V9�V���e�l`ޠ�����������Y=K=�'��֚�6�g�]z���/���,��(=��ؔ4~�M��_+��d?��#�r}��rrU��r��ٿ#�dG3�^��3���w�i�N��*�J�5{���Un~���(�޶Q�r��~4�ӫ8�����ɖ������ϕ��e�Ds�U��F��iY:�9O�'۸�����������;`e܆�R���k�7o��L�!:U�hՉ���[�y��AQ�,d��z���f��؇��G����x��>HѣXxjȷ7o��N>�.��4���U9�LV��c](WS���&�c�������%��0��D��T�����m��L)�]�t�glZd����ڗZT�*����YRR� a����,�v��t�G$�E���U�iD��b�N�Ld
z��}G�V0=V��z��yut�۾ ���H3��P�B�u�25��%ѧ(�7�N8�(;|�H�O;�ͩ�,�X�	)��򺽵d��i��)���/�ɸ	�g����.����K��J!�
���@B�L�1)W�Z��/&O��	&�#� ;���ȧ+ks���!��z��$�� �r����6���Y��/]e�[W�_I�"�sҕ�s�`G_�����l+4�`��hgkJ��W�E�%Z�����q�ƽ�%�s�p&&~���g���;ۗ����ؔcF�����ZzoX�����%�+��y��?����6{���i�1L��D4h�2W����?�?p\�am2��&i���
�\X�gkEG�k�*�]l��X<��<�,��=�z�y�[�q��+��Rɏ���:/��<�Y\[]eeRڨU�y���6�#�Xtp2�9���~��q��ڃ^&JRt>�}��?`��`�î�ڪY8�M���J�_�����J���݁5z����6l���u��9D��Y�Ҹ�8��K۔�4j�B��@)x�W���/w��}�m��8n�5X�k�3�����*�T�Q��䨉�8�OO;b�/����J��� �%�tY�͘���y�+���Z�=dJ�!��K��A��".�	��+y(=M 5/�Yn��z��@�$2����Վ&��x��]�p�� �mf���	�V����iJ"����R��L��*1�.��˒�ѓT���F5�N<z�mZWo/K�{SM���v����͚����䂣�a��X�A���������\�{���c���l�}�0wU���Y��k/<���(!�	�`#��j�_�����?v������o���䈡��៞{���v'i��e�� w��j��!��c�d�uρՅ�1��d� +���������K/���Q��H���y��wJ8���́���������Z����t�V:t��+���E��۠�j��`Hu�G�[����l� 87M�n=���eA;S8]B�z� �Q �c����K�]3VJ�bJ��R*�:Q
�ջ�g�m��u��n�
v�Do��`��V�Ǌm"�Ҙ&ce�5C�7���������X]S��@��F�e�f��\" +�&����*�fڧԦ�w:��#l���y6�r��C9{K��_y���_`��+���[jn<I��J��;$�b~��o"�x�I�	?|I1�OX�*��BNS�8S�H�Oo�i��w:��X��Z�%l��	��?IW@�&`�r`mA{�r0+D;�sM�!-�2T��%6��i���}�V,,Sk�R�ZgS��l���׬EjOW��ls�X͹}�":値Q40-S�9~��Zг��ѵV0���Q"Vu��d(�@��Jʶm^o[˶X�����}e�B��9V*tg]7.e>cON^��X�4?Z>�*CWl���\�=w%i��(���.^��3��Z�H��#���>�2��*�CҰ^B�b��;�G��>8@ƿ!���+��oV��|m��:��4�Z]��%O%�)'Y�qGٺ��z���Ci͆E'GTNX>.��c�U�^4H�@޻Ї�zD�E�����VьM��Ű�ܲ?��V"(w�B^�����j��F]�޽{{��%X��������$8c-Q)++���,���T�X�
�y)GL���?k���;�ht�@Ġ�] "k���W���l��o�O=�F��p��f	7dbx!t���4[��Ys�I�f����V� �جLx����2��Ƨ�,�?����K� Z�+�L�V��k�e�B�
�I
X�XU&볢	��Z-���X�Ԇ^�ћ�����2W��k��z2V���4$cX]��՟t�8��q�+_o'=ή�칖���a3�ϒ �iv�E�m��&��;7��rU�2
�\�I�f�4�@kԟ��R{�]e�abNY[ N[_W��k���!��*kdo���t�s�:`w��5 �6�L�k��Z�W[IiO���x��k���,�q�Vd�<����=�\��ܲj���og�^�H2�T`�������q�� V��c�1��W���Zj,�r�9�s-w��jVO��I�)]��`m���SҐY��ߦ�)�I_7u��X��^��2`�uD�����?�"�m��9~�d�>IM~�4>bR�Mse��9c��/�5�ذ �5kW�2�Q�K�Rp�G�b��Ӹ��G?��v�ձ3`�F�]3V�Z k�vS��Ӥ���+>igO�b���X���k\5lq�8s�*����!�"�E�	�P�>����)�ۋ���}/ʺ`�ܬ/���P���?��/�"YCI*0d��u�2������%��bpD\�"��� ��VJ���nN��q�V��v�(\���by͖6nH���W���&*�UJC�o�V����W��w�~�]��(��� ����
�>>��"���˒���P�-8�h/�u�t!s,d�W�(��VU3T�mt���&�s#��q���>l��{p1z����/�fL������GW�LԲT�H�v~���6U�Ҋ��!g~l��X���+`� �*��`wu[��8q����P
��1g]d-RH�k\� ��&] ��b�1O�&@!�lV�#_��=]��s;P���"���DC6a&��3VJ�QyiG�^{���
���Wg	Dp��$h����h;HO~��Ud��z�I�]~z���)C�8 ��yut���2֮=V�Z�*��1�ٮ����^l�7L�| �P�D��wZ�;��8p&?#���Xy 歴�y�h�;'<&?��q"�
X_�g�X�e:.`��(i�>��@�k�4����}��`8�
nW����^� 띞��R�Cm
�F���%��bU$ӬF�ߴ����6(�-��W�h�_��){���$����m�x/��{�N�#�u��z�-X�9"Lp��.,҆{�GkO&�����IGh    IDAT�U�NN��0����iܦ�le�A鳓�/r|��]�z���f���	'��k�QA�ܱ���`5 +=/.RlR�yծ�v,{����crR�'t+d���aK*I���֢��w���?�Ǥ�G&������UqG
�&"�I&�$��\�������(�������Q+X��3�j���z��W:��n�`��
ΐ�KVv������I������g��뜹��_=�q-y%b�+j�V0���uO����y{���R0+�ڨ�4OZcU����K��6���J�@HY�H
��c� ����B �='�j]�a�'�\u:_��r)�X�?�f���󤬶n�fi�V� t`�X#���"z2n��ޣ�m��u�/	Xk���%
�V���t=M������S�2��b�htq���6j�P+��LCu�͟1ז�+���ìUJp��Q����8���,+�~�]����.x�>���Ĵ+3�JR������5����{>�)0�Z��J�3����VoT��<S����sJm�Uƚ#>�l%j�zo������lU�Ɵ�ꩾ���u�ВqC(�S͒�>e��"/�{�~�.\��L���2#�R�����D1���E���9V)����CO:�2Gfm��sj�a����H�h��93���f_�������>D��'��M L��^m�n�o-��d�Q�?k�����<n��X�� k��7����؝� �ڂ 7x�`�V�3e����v�|���̸�Z)�v'�(w���mW��Z��c�H2Ɩ�-��F0젌�C�ʕ�ʐ�����8��`$i�I���,<	J�j�/!�8؊|�k�3�E�?�:��- @/8M��}�?�ڻ��@��B_YZ�̹z��8Fu(�я�^I)��� �����V�D%�֘�H�"��7(p��a^�U�m�la�r=�=�'pȈ6h�({l�|[-��|�k��^�-=�l��C	�7 ��I�W�<2Q��?!0o�
U����r��v�fH]�n��,��ɝ�tΞ���f֓��@�*w?a��[a���k�lW��m%zϺ.����|��*���T=�`����S?�鬽�4�ոͧ>�);�#lƌ��3�Y�1�`QD�MeS jCs�wdt^%�o���R�)�GN�Ȃ��e��$�7�C�K�=	a� Q����NɃ0-� 9<�ޓͧ�>�t�a���ԇ7�}1P���m���&�LW�z9�_#�r�����ֶ���9W:���˭r՛��b������n�m���qOI���"[!2/�� A�ĺ��z�Yg��	�^~�%{�7�U_��K���q"ҵYP^ړ��=��#۸`��^YȐ����4s��S�-	ѻgo�Wiӭ	�iö'��T��eʄ$��d/c$a�� ���#�2D>�&�y�;��`Ԙmѱ`��������;&%��A��Ǻʁu������RX}�r`e�&f��w���t|X��h�ȃ�������n��a6��*���ڃ�Ͷ�E&�^�/���l��3�Ҝ.��`���:�vh	37K��u���uR�CА��&z������X$�6��+ay)��UW0�t��6��bg_v��򘭷W_}U*O��I�V������%K���Y��Q��DM$�	������$�qْ��6�n)~��>�J�ť{�ǿw���c��c�
܆��տ���*+,]�ܶ�� ;���Z�,bj�[�D�5�T\\��+�jP�C�S)������l���a}z�����ڠ�k�%�u'J4�4a�D���G�1�[�:��f)��rj�,e�u������ho����j8� Z�JD�<Қ�ڗ5��A�z�����mVn��6ʹ��QP��*�/��ڭֻg�]!?֞Z4�C�k��%I��	ˌk��tow/�)�`M�Jf�С��JpE���_^���c�d��uD�?C#[��,GY�ǩhv!G �?Yb'�s2��,��6��,:�-�r����dU1��̱�r0�7���lT#�D�I��(þ��s�{@2U�_���*72�Ф���XKJ3Mc(�|!�p���ؤ�"�5*��8�*n(�r�6���A�*P��<Q�զE�j��&� �o���Խ'e��"�Z�AAc_�7�����z����cDy	Vp�2֟�r��k�U��B�$8`\�RvpMv���'�.���ֳW��X�
a"��o[��V��m��ʪk�%�.8�O|�����ݥaz�d��29N��\�_Z��:�l�|�/�"د�5H0�^/���` f4���}�c6�v��z\��ڣKXGIjٲ%����ց5S���w�}��@@��Z���v�Y�t"�z������������vV�X�;���mR{�1zK�e��K#$�ܤ��Bio�а��XO>Ǌ���=dz��Ղ6�ą�m�Q��KK����48%�U�A�<5���tCT�ل��'�9ۖk�)�}d՚�E�BG���֎Rb~P�^>����������l�jg���
Kzk�γ*-'5
 T��T�T��]&��A�{�)"����X�X��>y�/(��u����z��/�'L��z�ڕW|�Jz���т7��`�6���lh�h<�X@^��`n�y��m�
+8j��Ԥ����a�F֘�Ĭ$qNM�~�p���=9h� �h{m�,U?�	0s42�q�&��<�d�H3����t3��@��\g�{ڀy6�$�F�<�.q{�1r�q�%_�K#�u���VV�J�ҕW֊a[�D�_�(�k�%�5�M�Ei���$�ʼz�@?Wϡ� ="��Uv��#l�FmV�ܨ`�|-]I��Q��9V���v��:+X��ӛo�l�� �d��S<�U{��~E���.����R�'0�l�f[�t�m)��qW���*w�Ѵ�m�qR`��Oa$a���ĥ�uS��9�H;�khvg�:�OH5��{��^��UN�<_���\+�vD-r���^q����#V�!H^q�gm�*Ｓ����/5w\�* }���Vy������cd���3VV�T3z��g\�d�`��q���/l�:�����
�xGnC4�M�t�$�l�ݦ�M<�#�#���9���Wmq׃�?s��$3֯�n��7r�xӲJD�҅�֢=x�X;��cl��^vH�G�^h?��!����^���������I�@ ���š-ŝ��3�t:��L����R�E��B�=�$���.���眛7i��?M�~��\y�ȳ����k�g�S���v��H�X�8����J�,#lv�� �p�s�{�����z�"�ٲ��� c�n`%/&2Ҙ L2ܜ��	�^U!Hl��\��-��{xԒ�呦�+�_J�Ya�KfX.(E�yv�%�[*Rx��/\ �����S�;:�F#T^E�=VQ��)�{�cO>�,��>ǚ��ϱ
X٫��W���P��)�A�,��^՟�~B,Y3y��3R�������z�I��B,\'m�xq�:���#=��?��}zdc$A���ֆ[_�ÿ�JO���e���K�/�Rm��3�s[�d�W�])l��C�V�{�e"�i�o��`f��D����ۋ��e<G�u&�y5� �lX5�z۝�`��C}��M�¢���Т<2Q�o���!�K�������m!���0�� Y�!i�P2���sBw�R�T���-��u�����I���wvF&�x5���S��ۙ�M������ߵ秼n�8�հ��L-<��c!!p^*��>eM �fje1f�p��|�L�Ou�������=�٨��'�w-��b�Z�aN(���Z����+�Q=V�;��Aw�uxy}c��[���\�*`�
X������������U}��]�n��eV*`�dv�S`�GP�����_�k.����p˭�����V��?��u"#��d���Y,�y�	�;7î8��%�Ǉ�5��Ka@��;�A�H�T���?�A���|���=�����{%=���^\\a3gη勖Y֊8��qô�9�ry������x�&�U�c��֬�X�X	:�m̕���Tr�R��Z֋�w1U-gj.������يr�g��Ŏ���Z��{��e'�x��Ԛi���X%^�"yC=���XE����WǶ�50�@�C�ڧO�O�a�G�5	M��Z�	K�z�>�	��f��-��f����a�cC����Wt�#����[!�W��hF>��2��}�~Gk%�?_`o�k:k�J�E��_H�w�g�z���{��AD���W,� b9&��Ɋ���U#+��X��eQ��J��¸LU�{��]��^9�VP�2#���Y������*��k*m��Ex�3?�A�fW&��s�~�k����hW�ZSh�G���$Ha.nN�|������;��t�)�-/�}�3)�ݨ��̬�Z�����e6��}�Fy��<Q��mIY��&X#V��T�CkEy����/\��z�	m��9V��-S��8�����.aK��nok�}|�\�l9y���e��]�:`%�Z�HK��2t�������'^���\p�yv�Q�Xs��Z�Nf���UUW�f����S�3w����S���ɔ�+�+\���`��=�VE��Xx�5�"^�ixov�wc������,�}�����ܹ�l4���MVߕ�I�T����Z	|5�Zk�R����ݢF�IK�
N��욫���(t*xƬ���;P�5!r��	T��c���#�L�o'�p�������U�qւ�jP�j�U�*�������m�3���ƆW�*�{��;�x�ӏkA���E$e�;��C�7m��0b�	���m%�{�ձ�+c3]�ۄ�pI��]�1������;���l<(�����O�pJJ�Z��g�so}h� �4,��>���-��jO׾D�����x���[]1tI�nN�`����X�I����%���_+�`'�&��
7��K�iH�"��ֺ]�����ٖ�q��M�@���z���S��
I}B��Y:�TT`�^p&�F�����m�F�n�~�U�닯X������wwڛ�!`e��>Y2n#`U����%�Z�x�=L L����l�
։��S������]�x	*q��o�b=�ڛ_*m�?��T�/�Ǫ<VU���F�L���m\��Cy��ETv�%�l}9����=�A��V�	���Y��nc��o�k[���F�n?�����������"�P��ئp#���+������A�Yz�,�m�_ήJ�Ŀt��r�X`�WS�>Էhm���2?z���?/���.{������>�DIeC9C������T�����N�+��E|,��V�c}������X�تW̱��:n�T6�z�O��uk���J:�Y}ui�}~�(�D"����le���o�Z8�>�l�5���T��SŪq9/�Xw��������i�Uk"��Fk��^�$@��J�ء��%g�V#����-�àg,�w�δUkJ|����O���I�d�VjH�Jl�tP��O�a�z�g����l��C �����{�a���b3�[��$�SE%b
T�� �^d��n����u��V���������3t��������uP��Ļ�'QAfبA�m�ȡ6|P_�A������[ZF��oo�R�Xд��mX#w(Y��m�@uذav��߲�5���{�$2t�|��v啗�_�y�^y�}�`~������t"�{=�����W����=
O=��xA+��~�����?�R�:}��Gb��a,`m�g3�MT�e]]Yg_{��_X��~�X�.P�����{�^�3^�(I�����?�Tԝ��h�_~����׹]��Y��Qd��A���c���w�"��yy4	8���ly����<�ӣ	b��c���K9.��3J�}`[���F��e��.�-�����گ�n�͵���E�����d��v�~츣��|�\��?�ny�9�v�Զ���cM@��뮲5e� ��(|}�Q�:�X����
���.X��d��-�X= Y�s;���ḍ����n�4��Z��I�X��R4�+�Xw������ ��K	�X�Ni<V����N>l_���oـ� ��Qz{����Sm�
��&A>�6��e����P\�>����5��c\3���lJ�}���N��4fp�/?ؽ;g����Sh6�(�q�h��R��@����/X�Q4�U��V�5�F�%�ʞ�*
���57ݎ:p/�{�p*�\�,��u�-���w�r6��(ǐ��>_�(�������ڸR��b��6�Ae���>����g���3��D���pKb���l-���f���s��I%S��F3����&3PϚ�1��2rD7�V(�e;�U�AT�z��X�cmb�5��]���v���HXϽ�/�4��e*V��Ǫ�u{��H�$`�RO���$ܬ�u�5��#;³N9ڎ=lo{�O���5b����k*�c��۞za�=��K��KN`ee	��L���� *x���yZN!N&Y���.-U�@\�$xw5j�o�fs�Cm��I�eQ�n�4q7�ѵ�;�Ξ��Ԍ��O�FIP+�s7>8�C{z�H�	�� ^�T��x�*�m*��
������5�\���n�U}fv��I{�,$c����2��s��Tp�r�fl�ڹq���镬f�<2��j�kN���,t;U����, ԁ�ԸͰa#\ܮq;�A�8�<4T�@6��v�E6z`��w�N��/}hy�-+��~�/B�+�
a���m�wBp���r]�Z5\��7�ʌ�����d��2�.<{����S�&=������y]~'$�������t���X��4>���U�J,�R�J�t���*mha���'Wـ� ��烏�ۧ�Ͱe+V��Yc�L<4��5'@o�L����3A#m�����;C1���b2d�킷o&�3�ZT������m������W��鳭���L*V��"���:܈���G�UT0�`�ی:ā����5VU���o�b���d���}���ֲb��NӸ����o�ׯ��n�e/���:�o}=2������`�����(l�r�X�<�:r{Z.�ş��][8w��u�}N�v·���=Y]l?�ٿY���׿��ʪp�2MN���9v�%�!�.���>�E�n�e��\T���b�Wt���vw�� hw��	}���cO���M�7��]u��22ʸ��,v<K�7"9NG�����Eqi��/�__�Aă��s�L��hr��[��jVε,�j'2^�er�>���s��TO����S��(��!��g�%��M�-�R��ʲd���T8̲�'�Y��Π�V�M @�ͱ�0#U������D��K_��S��ӎ��`i��~��Y���OZ�4<�J��Tx�^��y *Ѧ|C[������xA�b�5�����J_v@����g��#{zC�������}<k�� B�5�u%,3�P��'x%=�8*� L$p^�R�U��5fL�`��IJ3�̺�a���خC3����.֧2��^�v��`y8���J�a�qh���0��*%P_oxtg���a!��?��£@��_kF�4�@����R{��7���_�~��21�+]���\�XE�G:��x�uڋY[�
���n`UH����c�S�ꩵ'9|��З��J�s�@CKi�A����T��E"��`Ul\3��~�9��y�:᯾�����v��D�K��*�R��.,,t��:$Εk֑oXc]x�=�$���a|��#�g���=k![_���cj�ٞ��b�S1?��{��OlϽ&�駝賦�j��C��Z����|�=<8ׁ�R��ʎ/2ڎv[N� �vb�y��x����9����N��Ԛs*��[\L��\��XaU��`��5̩ŉjb���A�K�:@����k��`�
NP^�z=��l(�KZ�y���߽J5��	�;Kvn�S�R�iX�C�;8�_�s���{�������d��yiG2����z�VYwlh��-��RV    IDAT`U5Ԇ�C���ѥ�پ�{��������?�g�1��T�"�)l�iEI�kPV���C�c���n�fP;i0+��K��X�V�9'�e��}�姢�兟|QڌW�1���3���c�4֎�E���4b���k&g����T��X5Ǫ̈́�U ߅�L:
۾�96�w�ҟVV��%�(�bZ�?%��6U���]yN�^�sV�@�D��F�'�
倧\�B���h�A�P�S�5	u�����m�@U�Έ�Lr_�E�C�y�	O��j�f�Z��k��F�US�c- �^=V�42nә�e�M��CoX=�\��PG�:q�Dߑ�Bs���#X�)V|���h(��%ݒe�m��9�h�l[WA�|�@����#��%2_�A�_G��������S�d�lY e|E�:D\7��(Qԋ��
@�rkr���M�o�Z��Zv��#4ˎ��kR�eg��Ygǒ׸/`�p�[�x>��ŸE�J�7��p�.vvh�:�uB<��.������nRk��x��V����~�a 8�H<EaMIŪ��U�`�vP��AJ�2 �{���=�#?|��&,JQҵ#`���vj��Lйz��DDM���5��;f)6v:/���W��eT�PK]���'�~y�����镩���p'I.�J+I&6z-�fݑ7m��@�$��P�,�Z�v~_]��5,�D���y A}y��/�_��r�<�~��٥��[���L�^Wϣu.��祽����V⼤�WQ���ߖ*�NrU�RGR�%e���ZW�"��Q.�*ÌTp���[(� f@���Cro����Մ$�IкԎ?P'o|uE�F@�YuL��s��/���b���:��UiDR��|,��6�/5�,�9�+���U�k���T�-y�:X��%�crs��dQ��2ڱb�2XǕgY=�{�5t^:���X��c��+�󷞳F�Γ:ߏ�Q,�zGօ��:�����S���-,\�t�:�p�Y���Y#n:����jr�I��qBӱ k�E�3�H�+�lgb6*b�	H}I�bLV���f�-�f{;�O��j�%ZDT�Tn���	�͝�A:u�U�hK�2�KQ��3൒�Ӻt�a^Xϐy2��� |#ϟ�a0o��5#7d[5��V�����Wp�~��?�c���V͊I��ߣ��z�s��z��~��ϱ�^3���#vDא,�d��*!G�DXe�-K���N�N7|�/��~<u*�TClh�؇8������	9��O�2��z�~gR����71E�m������+۰J�j��A5�nP�yڊ�'X�N�Y�Zj�[��v����g{�������?�c��$����6#��]��`]Q��7�2�p��m��X%^�J��*X�*і6�r��'wUr-.RL��푅x
1h:.}���ڒ/ʬ	�vY�*���mk8x�Kk�}�#V��X��d3�P��u�s]a��%lr4�UWj�^}�Z�WYc��6�����0i�����
���9`dѽ��g�C�蓩_z�f��z�u7���1�X�2O�c!�6��Q�*Vy�u
/7�����Q6jD�v�N6w��|�Ū���Wf�M8�4O)�B˞���R�i!�����NxU��=m	Y k+.*,�T��?�qrje�%3v]O�|E��*HI�c�v�y��PU6Zm(�Ӡ�v�Os�QC�W�b��ΚnP.�D̕X�1j�9?YTlN��E�8���p9?���**֫���l2��2�o����H�R��{��4�L�<>�[Lkn^�DD��b�摺\�H�`�c��FI��xzN�F�K��k� �SU;+�^�X[`���`����
�kp���K���ǔ�?�?��(U�rT���@�cM�)���`$ui�#Рl�U���]��vֈ귲�ּ�DU��%6� ����l�����`N����wZUZ
��]�Yx��b�N��i��88��Ĺi;�X#�%�;��#a��lP�^̰�Y&E�(�.�爰���)��V3�ו�����ZO띊�nur���:V��ݰC�0� @���*ܪ�)�m��=�]t�Ro6֎�����<T��;�{�w:�j���v k)a	����x�A!_F����7ޥ�5�F�W� +����5V�U�~��z�H��5�C��COi �p,��Wp��u,�5s����VT��5&��i��.�I�=�ħ�{�o��L*�l���C~v�q k�|2��2��(�WQ���|}��!]��K�u��Z������sO���:W"������T��|�g�[h~�i�R�/ȟ.���y&c��mJK�`�ݲ��$�`�ۈ
��f�Aĉ'`�����/�m���N7K@�
�Mͬ������ƌ�7�n�3?��a�vp��
����Xk:Y�v�XwT<��\_X��3���g����6�UkݒUܧ�����]-��<��`@Z�#T���,e�Fs��X֑ht/x�*Nt��9A�!K��;h\_f�/�����Ͼ��Z����Lz�����.`���Ͼ����R�X�I�Ѻ�ܚ��o�y)�F�%����.�R��o�^v�%g�(
f7��MH ���tQ�̬�8[�.��w?l_H�k�R�)�\
��X�޳�zm��g�7&���el�AK��
2	+]/��V�ZjT��bj�ٌ�&#xa��� [�̀*�4�E������=K�y�CN��_�$c1��S��ǺU`=��?�P�w���m����R�:���7�X��Xty�"������$J���g��\Ļp,�Kc�%)��ݵ�"5F��,L���~P�@�r �:S�H)�z��
��&��O�kU�
��]�r��8���1��.�@��MsHt ����
��X�o�n�H"���D%�P���,�e�05�/v`S��_�o�<�2Ե(�����Km���
.[WK���î�]F��Q��^=�����$��1���w`�@�򾚅�;�#j#�#��P�K
:�t_�~����K�$�U���5n�DϨC��Ίu��B�*�j�F��Y�n1_~�'�G���Jq�������O`��,=��}�%�t;Qͧ��t(N�I8���L��Lp���H2_��p/Wc����i���o�1���M��.'?��������{0�G[ˁ�w�>��/�Q��$�&_���nXei(��M�K֎�w�����ٰ���XʪP���༌+�����b�g��ߖ�T�͠T��w�X��Zt�u����� ����X�d��\�:䅙4��V�ӭ�T�9��^���j��V��X�t ���\N���\/��1�V_O==4̂~��G �n'������y�5xqS`��R��WX�g���5�cM�
.�9I�z_��E�F��MC��HÃm�o�١�Eu�}�e�B��s�U�Qe"LR/���R��&v�K`���[:��>�8vQ9\!��:w�XVvF�յ�)Dˢgy]1�ݴ���Pt�k���mֆbLB|�R2�g��v���>���EJ�"���+���޷�_T���N��2$�`��뮳u��ߍ�Rbn�k�!6 �z��Q�bNLb�//C�O��h��˗ۛ���}cVvdLbt�h��[x�I9x��G�͗A
�����9=Q'{�Uy��JFRx���T��vMD�g����ZRP�Cm*=V-�q�bC���uT��	#�O������Hn��	�t�2����$��詖ą�8����;�AU��^1�df��0hG(�f�c�T���N;��?j�E���G�D�����.��:e�&�֔ ��w��2+��	�i�,���'�k�i�M,�j�FT��]�v�Nf$uY����F�agϼl<w�؁��1V(��*
�f.�;H�b�7]y�����X�3���8*`�ǥ�irϫjE��������UUwkq�ym<��U�N��,+W�k]�Kr�S�G㈢�x���X�ώW�I�
�酔�:�l��Xw�<���sA^�nAl��@��{O���Ҳ��s����BYc�!�Xu ��h�&p�I�Zu�[�[���	�5;�o����Z ��u�~^El�j��*D�Jj�'p�ĉ/*ƄU�!3G����o��pJ�O��r���dUxl#ʠC~�>��E���C�©z�2�~�(�+%JG�܎�vEI�1�_�Au�F�+R9a�b�T�;�N7�����5�Cv��P�j�`��Vg[M
�}��y�$ͽ!�O X�cܦ����L+�`�(�m˂�N�XjU+�c���Gn�]H�yQ�"n�v�7o���	�2}~M>�>���>b�%dP��QG�T�n�(�\�%%
��B��=Ľ�wR�;�u����'�i3i����p���Ϧ�,j+-��4W��4��O=��<y_&�W���g_~�^�Ϸ����V6���"t&��p�߷�$,���,�w�bT&�j�sR�>��3�N<�h;��q�>�Ҳ�����}�ޛ��r4Vȳ��Mq�-��4}!s�U��4�,���6E$����=m�vr��Hv��N&$/I��cj^ͱ��^�J��X��K���e$kO�?��u'\d3��E����8$�c��`i?�n�OEL)\FM[��u�Ì�!%� ��ӽ�>s
kYTp��7�;/�'4�!F1�,h�QB��p�P���!�� =�����k'�ie�H�$�����+���"��:���Q�F��|,;艧�f�s�uҞlb�W�>wd%U�	������?R��jߠb�C�zĵx��)��/�߽�;6~�x���٣HT���ǆ�G�q4>���7�JR}υ+�`��1��z�eXi +�!n��+���iSC�e�e�.'����C�%i�@��_�2���G�S^���Et�S5�рs�fAc��kp񉦎c7W��f���!��Ο��:���n�M_`o���}6}���2H�H���Ύ>U�.�$~0�,�kQ��|'>Ʃ(�}`�!@9�tk\�R�X/��r���t����z�=���6q�J�q�h��ݪ�'�w�qa Ω�f��a{Z���4n�9VU�;�mv�kc{>��r�y�M �Ӧ}ė�����uU�'n])��l��s�)v�1�a��X+ļť��[�۴yK��1O-#!YT���i�\�����&����F3)Jzr?+��P6������j����'�>_`�y=��H>���yT�k�V���VW�aA�Z(�zs��t�������p����T�GY6f��[s������y'M`��"�~�Ï��^�`���c��{�a�E����D��Tʪ.��T���aR�����%͠{_5�йiD�,���!^Y���z��&�. j�sԘ��U�l�uVR5�Q�*�Aؽօ�v&��J�1�s��j���G��7�no���.n��+����1k�\�p(�s �B�x���wB�� X9����J� X�Y`� X_(oRŊ�g;+�3N;�-�-[f3�+��Ѿ�-��{��!�S�6ْ��J�q�m�#�e��X�[�9���Jjc�3ۆ�c���`?������;�WWY_�mà
�1fݳp�B[WV��@�mBm����TF����ZX�O�h�K�#�ڲ��퐉���N�~�,�~ӕ���̳2�-2�T���	7���g�Y}>����D�Эvv���U�&e���bK�z�eW���n���_`o��Q@��H���l��m�:�O�3��M7��[��t�kH�O?���˓B��E��*6N�Ɲ�6�t��}Û���U�j�@�����0�ѹv�9�P��bA�߄�v����^ռgp�k�Y_�d�������*0 (#�S@�|W_�CC�L�<L�.�J<����!���� �'����0��x�\�%��3�-�Z��
�։�� ��&����k�ũ`��V�$=�L�֪u�#?��<�����V����Uk��Yg-�¾� � q�iZ��J	��zWŮ���#9��a,��`��&ёҦT-{Z����e�H���������l��Ly�$ѻ����𷕮d��Q���
5�.!Zt�p,+�~l/��b�hv��E����*`�{ϣ%�Nk����\r���0��7������>���N��ͱ�]Śq��7=_ސDź��z���yŪV����0�����$��f�sѝ�]��AígQ?��-��V����3n��նq��;P�Lfv�]���3*��Kk�λ��:��,I$��Y�O�=����4����@2���so�G�~�j>Q��3$���m^�h�X�?6I�.*F4�Y�ώn��d���T.�8���iMH0�����vۃOc��*�X��B`� ��P�+�yƁ������\>��b�����
#6\��
����b���F|�a�9����j�FT��U��;�m�Q|��}2�� a��q��<�S�	����P�60�Hs��Av�1G�i��z�c�[n�.-���mg�yN�ë��]���,��zK��f�\��{���g3�����Rfڳ�{Z+=ZQ�)u�=�2��7���ST��<W���3���*�Yv��X�E���,��j9/u���xxg;5rBK�[l(_K-�{*�Q��d��>��
�>,��O[lO���UR'�@�ki&�u_���p��Xxm�@5�� ˺�֚>����m"ny�,�Z%�j�.�Q�f�+ҴD(Յ6�sұ��d��/��/<��vι߶�cv�9sfٽ�����^^��7�/��{�{Ʌ>��Y0�+ִ��m��g}`=�ڛ�+mJ<�� �y����J���owC�X u�
�5v�U��a�,�����\>���>��l��,�����$�׊�g߉#�ΰi��Bq�M~�%R'>c�4�5�ۨQd�[��bv8�%ؿ��O����|�+0]#��8p)\څ��<6B�{�J�ᤏ�����;��xxu�9]��0�r����Y���{���Nb���,E��1mT��>J��s����f�*�P0��̛�T��]�};p"��;�Ç���G7�(Gy�W��i���;��s�w���+8�h��ΊuG�2��%�	�`��B���L�XFP����|F��q��"������ �We�|W ���%AN����ZUDFj�]	!�lu�͘3�>�1��s ��������w9��,�FPĤ���>�`���EL"m!�`��n,�ΔxI���X����G^�u�׆�U��kv �Ҵk2	:��?�2�m~{�d[�p`*1O�m�f�"�}D������E�TMVH���B�MN��>���c}����ӣM�&�G�gw��<o�
69>k�c����@}،D*^*�/�e,��s�;ӆl��ϵ0�W���h7P���7}��9b���������T�V+֯
�{챇���y���$�S;l��� ��Z4�Y(�՗ϱ�r�2 �#N���"^�d���ʏx1.K���o����/������jI]HՌY}-�O�5/�|E.F�^y�5���翼�J�jKB��.5�wo\>A{�{�5/�'	���<�����q��Q0'�����D��Ui}]	��{[Gb�[D}h4FC�P�^�=�Fz����`U�Q�5�X�]|��$�P��s�9��.XFNb�۱Sܑ��nN�ۈ
>���g[�̝e�<��ϱ�ǚ=`�%��Ӹ�;��w�c۟M@���Ճ�c�KR���F
S�,	l�>��l�йm��� F�U�ܐ��P�YQA.V����iK6� �xw3� �z��Z���	)Eӱjm�-_SfŬA5�u�+C4����� Yl��{-
��qX�(�ݰA�{�����T��k��bxVU��(��-	��^�� �k0�b��q�t���O0GK��V�e	���8�5�L��{5'�QC>��%�8dU�~�������:���U�湦��8�C�7�e�?�����s��[�+��MGb�,�re�?�'��yVQ�߻�<�xй����f�*V�1
Y��u��E��F}#Tp�����\���    IDATYC��_�b=��sl�=�t���܈
�D'%�:�C������ng��9V]	߀kOT���X;�v��ve�_u�M��{���H�9�N9��ݟ��[&A����r5d :��n�0
�n<��zo�=��S>��I���)L8�����)8�F�����y�h�)���:�?��*8����b��kk���	�)&^_��T+�p'@�+����qmR�z�}[2b����ָx�~��{��������U�
Xw�5rb�6g/E�`	��x�5{�ŗ�+Xs�C��k����mώ�[�X�.9�Fd��4��#~��/������>�F�`���fg37OKM��$��Dk�r��EfI�д�]#|���z�����r2Ru&�&%4��"�6�
4ߋظb�K�X��4J��
P�aS*xS`����g�+����0�V�6)b�����o�&J�g����d�h�/��[8.qz�:Fz�CB��ȣ�uJV�!���<ԃ�׭#|%�j�O�8e���ճ�����7/lh�|s}b-0O��ZBR@'�v�Ře;�q�j�fr�о����~��-��z�E��0Ж+V}F=��Q#�
����`�b(t�~豎=J��m���V�~%`=��gzl�ҥKMA�����iD�Q5;��^}��.�Ծ�x"�b����-��0(^@�����oE=s�[nF�$�ɷ����
\n?��+C�/�.�U�m��=v�s�=Պ�V�-���!���lDڝ���Zi��w��C�O?z����E�0�8{��S��*{
.�2h�/j��\aKV����C5�uX&��řIh��p�0���]�5V�x�ɏlXU�4���ͣ]���
�ʑF0.ԅ	����n�(>N׎r5�rТW]Si�����e�M����q�*b�v�|el�g�º�*8/i���Kb�0.N40�-Orm�%��� X��|E�|��/��sP�k��{�A��aX���PK�G^n�1yY��LH�:�iP�U?RB�wD��`]��a"��F?����nM�
lZX��� dZ藦1����P���t��W)�1�|$��8�B��D;��C�	��y����3��瞳��J,����~kXE�~��MNtaG]���X;��m�`����'Z�3��6�A��\�W�ւ�$�l,������H��\�zŕ�x�:k�VU����o�Ǫ�4v�шcX��X��T�u���y3�b�XSHc�xIT�*V���P�ƎHD�ƦB&=�0zE�T��;}�k`a��"豖1`�5u���_��R��h_�٭�=��Ks��Gm��5R85d
��1Gi�?u�{��Ǳ��Ҁ"�I�x���)�u� �ɲ"㢑��'M��w��(z��<lW�}]���"����-�70k�Zd��o�Q�����n�'ݦ�n��J>K��El��`�=�؝e�����.{l\�V���{�����Z�!���Z��SUF���d�0I��b4T�2�����a2"`M�jS0�N���+d�Q�<�K�8�!�ﺫ������a}��(X	[\$sG��'��l���>AT��H'kFZ ��w ��_Ȃ)[Y�3�#2�צ>I�ߧ*Vx<m-%�(P�)a�1�_��qy+�e{�K��c+V76P�+k���z��ȏ��T
�p���	��K�g��^c�R��5b���b�1{�{ꉇm���o�׮�^z�i�}�=��k���S- L�O�%e0o�ԉ8��7~�����_���f.`�?uE8"���X�1�w`%�^��E߿�{��gϴ��~�3e7�X7 k�B*��w�দ6/�f1��tf�5C+r ��T�b(����6��:^y�H�O$��mXu�D���"DO�0�G��RkpQO�vyѿu��d���h���T����~Ǟj]�i��p�}���S/�
��	M�N�^=�`�>�X{�å��#�;�ѷ��u��6f�@��G�>�nU�id�%$s�P�i�;!l����8�
���ld�i�`;h��>r������#)��F�;�PޡC�}�Z�,��קۣϿfm�۸��8�P*���]M�B�ݣظp�&����cM������D��$`͡���!`�Q��zՌ6u��5�]�b�T���XH� ��*�wY���)g.�ۨ7�Xw�Kd��-I�&�z�,��#G��Em'8(��D���<���L0��h!�lPՒ5�UNc��3M1a\|���G?�_��"`��&_=O������ЯT��jmR�K*#�p��D������ek�r����/mX5ʣ�p	z��hӨ�Ҹ��ٝ�v�O�޻6'�|��c�-�����Ç�i��hO>�(��Y3ӭ�>v�	' � &�i6�7]4&��B�}'/�Tc����ء������E��ǟ&P7������
�,_m�Oy�:�X���������#�8�����W�-���9Ǎ�i8�H��-Z�g��9�]�<�����K:3&)��[⼔�o��t�9V�ߢ���Ŧ*��OXT@ۿ_/޿�j#��S�&��Ǟl����|�w��f�]?��7����%�5����<h���wXyi������6{���h��ݷ�,'����E�l��eЃ��̱%��O#<2��#^
�9��T%3�Mw���?nX��ח��ϗ�o~#� ;��c�C�����<������С/p����j�v^�k�W�=>�균-��..��k�v������SP�����=���N�qk�#ա����s:��Y�P������֑��vÓ�vZ��"k$^jR�7w=�k��fϜe=z���X�hS��8�&�`�&�f�ÂA (���E��UoL��o,5S�����~�j�U��� U/����,A���襆�E�#hw�2��9�}�~Ec':�,ֆ9�M�m�T��sW엀Q�]�3P���n��ц$
�hU$�<ʃ�9��HN��[���L.UhY��@��8�e�Ӈ�>�L�o݄�j����*0ڨ�����aL�/<՞yy�=���--�șFm��p`U��*Z��X)v$^����ڈa�m���v�m��K7�n�b�y�e�(+��Áu��YP��#��ǟ��V5�U-� o�˦��g2�P&����>��{_:���.�MDf��nO��KO���Ҋ�W�L/�"�x�	�@��`v����ʫ��
/�LA����:q&�N�أ���{����v�I'8� 9wA����$�����.c*}:�K5��KT��զ�{츍�޸ ��
'����k����r��l���֋JY=��|��1Ӯ괿������'xc���/v/�8���믷5�/݃	�BwX�;u��`e-��e����CNU�����Һ�wp�%���VӍ�?VWzr3z
�Ga�YbӤk�m��P6*"���;����U��mF�Xg�dc�NfN���`J��\�Y��yTfX%���o*G��K�$p��2H�Q�tjп���o�Q��T�j�/��~����Vէ~��K���KYҮ����ի����,��+W�O$:|��`m�Z��OhaS�k�t娊�gM��c4����(N�~&+�_(��b��Xˤ��P��=���Fn$ĒHJ6��N=p�EQ�51�W��v�kӧ��G�~��4^AOP��[R����i�b�>E=����,*x@��<b�Gu�<Ⴢiӊ5,�ؔh#0�_"G�}�u!��M��و�Fv�vk���)��zÉ�MG���3M
W*�Y�h�T�Xl�9g���%�Zt #��H��w#@�����lղEx�b	��$��a��}�Iֆ�<�@;������Ȯ%
Je���Ҫ�z�R�����f�����zAxS_�H�+��/eg'�wV5���������-�K��v`�8zp?;h�8��%��Б�����Z�d�-\��Y���eW�����d���􄨂Ac�`-�){'Tp;�Xe���|��8 �8.R��T��BkK SkU������`�S��a�lZ1T��3��D�q �\���p�K��㖆;�X��t���a2�?�M���~���6� U)#~��tj6T�-N��^}����u�_yt�t��%!��z�kҁUԮ<�]�V���C`��Ń�Hf�0�ϸHJ�z�G��x��~F0�P�t��£�%E3���5*V/��L���F�XԱuDu��[��EK�� %*�@�����hC9��d��,�U �hW��r,�Qh���>����F�L�У �ɍ��f��s!�;����q����αH
G6e��I�o�d�����X�[.$9/�(��&�&=��m=��:���U��a/.^��%y'�b�w�?Xu~#ᑀU�%�%��v���:͆c%Q��:���zc�Tyt7�9K�"��2؅���^}�ȪX���%�`�dǡ��6*��F���}��O��1k���\<+EUh����
����H�^5���x� =OQ(�;�]�#賺ݯ����E]�Z[�����I��I��R��
�h�"[���.��jp$���g��ŸM�.Fޣn�4�p k<�6��@�Z k
U�_���"�X��#JF��D.��E�,�'\�+����E*V?��<��+VUHt���]ԃeL�K�$�ͱʄg�����X}ïjP:��\�v;�g�-^��M��^��O�R����o�28X x�&�z�]����CKB�:������H��C�\�^��.ö<˃u���Bf+�s 4J�������W��}%лm�xf��?¾}��n��S�̹���3/2X���.j����X��?Y�Y���*^t��u�pPzݣ����X!�S�4S�K�X_�ku-����w�.�ICc�����}�����4��U{�*�1`�+�WaO����3�S�e���u`Uu��S-`�1c�����V�(�/}�5V7]��*`���KV��3�?��`{�O8T�}���L~��-t�$6��a��>���Uµ�1�o�y���Y��QV�
`m�f�%���(�I�D�-O*F|��o[��ur[���{�$AFԄ�d2��5qҵ���G�S��&X�� B�M�̪L�t�����l�i�`Ƨ$Ԕ[Uk
ߺ �<έ��.�8�d[�-�Usrɸz,���\�x����$6.)'�{����
�	ْ�r+��"���c������.MSo��*xG�cuZ,d<�M��7Qd�!��Z����|��Yt�j�FA�22�i����/iï렎Mx>�-/�Gx�Jiw2�����3^�H�yUI��B�u!��c=���u�R{^�J��Jp��VBI0 ����fU�\H��b�2�3̆�Tp�\��`�f��ޗ��%��:#1��>��uK�-�XEc7kn����N�YsS�/aYN��=��^v�Co�Lc4�`�n�w���QB"Oݛ��[S[�Q�n�{.�rS�
_E�u2"�ߩ�ߣ62�RLZ�(�7"���N&�:�R��������0��;������Vr���D��t�z��$�X�'�)�CM�=h�?�
�XӘ���.��w+�j ��!�R�.��b���7'fr*6ht2�m���G�d����KJ='��Q2�gΰ kT�,I �V΀��@Y�(Ar�����G�D�N�]���lE��.J=��r��~�/�,#B`�}�b�h��z�J��I!ycjM�j��C����xd�"O�T]$ kR[���+ �**�G,)��qy�&��q�X3�ڝn��%��W�L��ϟo��Q5����"���]��R️X��Ed��PJC�C-�}�����w^�	�ǪqV�����^ Ɗ��Ϻ�����S~*�N����(��F�h���z��+�hժ�S�����s%yDE�<nY�}3��������h������с�6E���F̔���j�*�[ց�����~�s��weU��/��j��TE��&=k����f��} �ʦb�$^�j�+���}z�]�7��!�,_�&�b���R}�jOi�`��Ů��J;���������b�xq�Q�ө�z�TS�L,T�{yP4�(����ԏ��~N}Y����:7����ԻգI�~~&V}ݫ|�X��YۨXg=?�U��+OU�CϿ�}��oX������ ���V @T𸣥
.�m���͍��Jo��?����F*�6�+��*�~�t�D�vt� q�����"v6�V���*Zw=a��ՙ	�[�@�=�~6��-�9�l���Eԇ�+� RP'3C+ʶA!��{/�^�@R�ޕ�� *���U�N�۫A��!�P2rUր�&\����G.*�`dmVSUfN��N8hK��K��7���6	 WW=3�j�?Y�=5�]��3��吒�E�R���U��j�.*�x�6��$ʛ�M�]a5+�X\C����W\�N5םP�z�����.3���������O�T�ގl]n0|��7��9Vx=_w֢S��ILUz4��u���'����#���?�oN�Qk֖2�xIT�*V�Π�s��o��@Uw}ж	[:��K ���� �u)�� �o�6�&b1��J���"(U���@�Nz9�:�d���V�zڈ���K�����S�V7(�}�&�a{�A���)���΂�Yüm�"R&�MU�\��̟��+8k@���ܗ��S|" :�x�Ӥ�z\�k�s��Sh�-���|Ԗ�#�:���t���T8�+foC�,�R���G�@��t�Ţv��6S�*VN`��*M���=�5�����o �r�J�]P+��9�<��6��;��zC�h)�����m\��́�,��H'�?�q�o����v�#�>�:g�s�_X#JWբ�`U��&a*9a���ih_�f��tp:���LY�����������Bä��Ül�FX3J�$�J'%>��E� �����j'E�?�&|��aR�2��Qרp�D
FѾp�ԃi��VCStќM�B���M��F��ˍ����T`�E9�f��8(޳O>�.<e"I��w��*Qm��o�̩n�U����zQ2�ssJ�*����r��l-$w2k���8U��5 �R5��%_��EV��y�C�1�E�6�`V��#��mj��h�Q[D�G`�N�ѹu�e�0�<oЋ
Íc�z�otߌ޿���/��X��*������*͚����4�	�_�h�����܀]ڠ��.C�5��%ϊz��#e��齨a���E����Ъ���TYx}��)~�`���6}_��k����ts��F��� XQ���X+=��z���c��5Rn&"��"��K�n&���T��&�a��,#��^{c�My�m[KXHEJ���:=�\���G>��U��؃w�m�g@��z���� ������i��>c�D�:�ޓ��H��i�NU��^�Ht˜G=֙�=����"���L�ɜ3��D�K���K[P;X�q����U�V����"5s�H��'Y�fi�(��}X�'��׶� �Kk��VU�V���}���b��BF[
<�G}
=bY?آ`��'5iav�.�%X"������]?ɒ�"�&�����&���R�ec�� �M��[1k�a�MF�7�i�TJ���ŬP�ͳQ��~��q�=�C��*�M�d������s�av������3�|��$Do��	*�T8�Qg,/��f�u#x텼�̸�;/1�ZLx�=�?��ڝm	X��%����ﾇ	���y�|m[��UL�;����Ǝ~6ꇨ򏨛����D��{��X�y~��D�hW��VW���j��w�~���U7�'S?��h�&�X%^�Y�n����y	�I���v���HFA-�b�D��RR/�����'k��>�6��'��� �;)�H�񕏠�:ԥt�@�E��֞;jkE���
ʺ�I��A���[ﰌ�~n�/5�*r�;R�_]�����N;�(�l��3�?���ɸ�ţ_�d�Z+�(��T�*<����?�}���Xռ#Oi�    IDAT�����AϚ�����f���攡��0�b 9o*o"L�#��b�Ӫ��u&^��m5�G�u���!�j@�ҁ5�p��cK��A� hi��.��
��g(A�g|}`=�ڛ�VޔxD�	����A�4UW�]x�y>c5c�{뭷|��W��i�`�
�rhVJ��+�/f:Xy���$��%�D?��:����D?vw<(gx�Y�3JX�Φ��{�=l�޻#���R#4b1���}�Cfq��G������@ވ�	z���ͣ�EG�ң�_��,փ���>�g���K�^�O���%� ٮ�c�2U�.x]�IR%���\ϸͪ��w�~h�%`����n�_�b�@):~��#*X7��B݌�o��M�U?��n���[�vW��� ���+/=ݛ�M+V���>��b�f�ۥ�b�	�_���3��+Lݨ@�m@�z��ni��"G�m~��N#���)T�AkӪ8Im}���u}���M&�)�i���*�K<1���ݧ�LѶ�Ukp�%���c��U��w3czCH�I���K���Dزv�-u���N�˾s������je.Y��f.Xa�ix��eiB0��B��"��\cK���7(�71�m�/��2i�%'V2A�.l�T@ɁI�+PU���gêW�*�b#�b���V;�� ��_q���O>��g݃^���X�""C�Co��G��{�`M�;�Ӿ�j��K�H��nJw���c���O�����Pk9��h�fY��<�5����ѷ���?`m!�f.�K�I�G�jɃv�:z���.����A���+l@�x� �~���v�́6S��S=�}�YgټY���s~A��EZ²����_��� Z�������kw�$�buQ��!	��P[+ e@��V؅����NߟJt����ɖ����;��q쨒�$��=�����>G���E|�6����n��̌��V�_X����"�� /����j���8�{]������ -B������ ��:��ݔ
v��RT�N`�&��?�s8�*�I�� ���	�B<_��^�!LQ�U�ߨm����6�z�ĥ	16�&��A�*�'׳n��jg��l[T�����[��r�Ϯ��K"��=P����+|��N�KY�v�����Y����uK#i�-5��]6a�h;���E�qC��_]by�y7`I��l�X��G�'�;��{(Gs�9���x
�@���R;ƀ⨺�׌J�N�r�sS�� �ke�b�(VT������d�ܝ�d�߯O_7������)UIB:L[��#���{����-0w!�qM0���=����s�A�5��֩��%3X�9�L�{�mQ@��z�W�ni�c�VE.�	:�C��I�?|A�s	�%6�=�X���z�X��4V��:�;d�}�O=�G����ԙ��cOX&qA���dn1��麚R@������\m�����?�����[(�VE2�G�I�-���aе��JT��եv��=mo��+�o�^m��5�H��˅�,*�Y�F�G��s�J��D�&�cMjETc��]�L�(*8Xc�/��t!���r�fѽ~A�4l���EJ� ��H./�%b_�B��v-[��M{���O?�I݃�O���F-�j�І�^@ENI��⏊>�Mt3t�j����K�m#�z�.��i�$��Qv�*s�?|la�\o8E�$-�
{�[:��VQ|��f��K���X/c=���=��[k��<��(�$��V�Xm$ja�/�ؼ�,2��q�ͨ�L��+�=rS"M%�ɛ)"�����˿�n �H�*�ς6�3�q �ч��������,)i����b�L���{.�7P��9hLI�h�|����6�%*��R�QWlܨ#=����f>�n��%��
��3ޙ��pѷ�)���v췿!`m�?�=>Eۨ�y�-k������w�ۨb�����H%ы�G�b�'�ֆ�B+gF+>���?�ظ�#�*8������]m��ϱ;��g��O~b���㿬��Wkg
�g���4`oկ�z�VAn�I���5���3��'�����QOHAݥ��K���#�m�)��0�����}���l�\2@_c����ʍ��e���K%��5	��
v�M]ǆ1���k�r��H܄��(^���� ���|aL����PlDVD�FT���O��tsI�'���F��WH9��cK�%}=��)^�:G���w=�&d�X
b��a5�R�O~��2�� �#.�j</EL�V�������E˭�'R�������@(�
�B��;R�����^��ܛ+jxQ��� �6*�;ﾟ�{��% 8՘K��l��񠍥���6��+ڐ�1_��0��sq�K3�)�^�&1��&�����i�Y�<Z_ҨL���K����<x��=w�T6�ծ�9���G�|����0�Y�h��O9�)}'X�1i�bu`�-!��Ѓ��C�:�� _��T�#��T�ƌ���g�A���`w4���Hź`��4lX:3�4X��w_v	�M�R;Py�H�# �ku8b�h|0�(�X�-�G��<֌�6��S,e�Tl�P �>� ;��#�W���-�;�=����P��g�<����8b���
;����C�#��޵�v�-w��
��Y�T��l����`�I�C���n VU���ȦK��=KT���,D����siJ�{qC��K�#k�"J-�FY��l�*�_Mk�*�
W��&J5ݼ����˯���m���k4n#�3���n�Xկ��c�ONFz�nG�B�׶t�+�R;Q���X�o�����}����Xa�hj��h�U�-��{�cO=�W����:��?���U�7�ICj�}�D�jщ�^�.'q���q���=��t�ϲjT.5�V�{x�闭�����T�ʗVT�^AUY�z(ʙ)��C��!��{ V�΄�U��n
E� kJ�믹�B����>K'�[IY��d�����'x��'j��[K#�:PI3��ql����^f�T�z��x�vz�g3�fs�y׉nX�k�ڏE(^RA'6���t�Cևb=O<�d������`M���4�9U����Ϲ��M ^���f5�o/r�`Q��'�x���j���R�WcF�C��4/�������#��鹲���c�KQ�����XC*��s��<ֵ���y��c�dwV
�F"-��c�ӧ¤v�5w�}J�G�t�e�*4Y�����N����HQH���=��v������]8����z�ȶhٴdvE���n�><���ϛ�#k�M7p�i��{��n�h��E��PE�D��\��k+�0#�N>�0;`��\������}W��3���^z��@?�O��T����J��_ZVaw������A�$��8Y%�Tα�!o0���s/��Y�b�͙��-ٲ3I{�� |�[�#*X�?9ЦG��Εfy��#�E*���B���~ֶ��m�v��#�Ԣ�"�g�}�&�?������Wp{Z�;/E�qRj������@N���2(p!b��vQv2�[���va'y�Q��J�5?�9��L<��z�JWV4�C{ժ��d�&X�q���FoD�-#ͻo�
�qT�:�V�3��X`��ܭ(|H|j��lj�X�ۏ�?�*p�}�'me�j(�J�c
�=f����&����v+��T�ٱ'b��\c���0�m2x��=T=��b*D}?�4��h8�iA�Q�x��QUU�]v�e�������>�f	��7���'�����A�tN���6��GX|+�Ǫ�u����*����m�ޣz΢�sa6��J��k��o�b� X��e���s���c�j���cSA��-��8�h���ع��"1��>n��AdW�^���p��F���<j��à,
���)����~�^{�S+$�S��4�̌6YMe�x��#.�?N�f/��������0�y3#=�܈����V�
�^,j�|�ҳO����'���U̓�Vc�R	p��i�W��<k��^��!�
�D@K�7�������M�u����C��)Uˬa��Utub�pVV�f	���vP��%�][zD,���ޢ��H���pS��u�F;�<<N��\}��~7�7�J;R/�]9.5i�G�q���b�m��7q��O?�[j��F��DY�q���l�5��=��IG�m��/��4@]YY��mgs�R���0G��X�]i�=�E�ڲv;�ye���ԛ�Ћ��Z��)�,�C`���V*�?�~�g�����~d��w�9h`֖ukڈ�\���� sѢ��dذ!�m����&�h�cO�ao2e!��8z��떁U�=�g�^f��JU�~Q�b��A�&�l2����퀃���߱7I,K���qEmp?B`�T���Xg��4����u�g{l��U�i-��ј���X�X{�*�q��s��C�F_�
�8�ڛ�+mJ<��T�g~�t����s-ر��M�|b/�aC�Z��E��6w�2h>MV���c�6�+��ʫ|G���2��ƨZ-/#Ѯ��J����M�,�޽{ۚ�� A "����������[o�f�Zh����"�%qI�*����F7�S�܌)����nv�'8�׷g�{SgY&�,Frf������*������__�.(��E,'�񵼑�U�z��XEGG����=jZ&2�Pv�n�^}z[���>Ĭ��"�}�`����G]�
�w砤�ʏX#ձ$��Z�.2�y뫾@�~xl!�-���v��[�k�#ZKIϳrf�rQ�X+Z��D��E�㝱q_��_�=����t�p������XrS�}/[i�6Ҏ9`��IJ��3V�B�-�<�-�h4��Z��'_��&,Z�<"�VP�-���X��*8V��w���@�Tm�>�k�I��^�w���i��A'����X8iY�V��l��U�ћ�/EPĴ�צT���i�xi����c�w�#�_NW ��֨�4;���)���ɧ߰O�ᑀ7A�U~�X}�_S�E
���R,�{�"
1�xI�T�걪E���U�2��������x�U�:g�B�c���K_	XE+�U=���۲��w� n��hp�����ܯO/�1w���RI��=9ƒ��ڰ�c�����cV�1�(<�\k%զ�� 4�;e�����uuv�5� D-V]^�I^^���g/L�ܦ����hY�/쒜b����D�7p$ˎ�&�4� �����sO�s��H�������b-I9����<�
��r�]q޷���W>Zf��1k���`g'�Tk���/�
v�wc�Va1��Z�܁5��^������X?fg1BD�X��(r)�ފ5��hW�4�y9E��}��3��E5��S~d:QR.܊9�_�%�9j�z�p�9�����+;9�-PW������1lOK*�g�m�RȧY��N`�*������������D<���F�zz�ٮ�{ٰ�H{(�ͨt	Il��&O"�6�6�y��δ��+lު[����Oܗ�7#A�|��9`�sS �r@�Te|1p^��uwޅ�aZbؒ��S�����
��e���A�l��A��� �h1 }�aD�Ś2[�t��+EG�)��8����8����� bc`툌�Xw��M�ec�XKo���#��N�������$�����Ć!��ڨ��k����e�4�g���؁U���9sf9�6��72�؂xIm_y8�?D�5c���7Bq�Mϗ7$�e*V��&N�h.���+�H=�>���1]|>C��
� ?�����󀳳�����k&����B(��� ����(`��W��ދx��� @@�
B-tH#	��@H��{��k?�3s2�L �#��G�d��9�y��}��k����/�緼޶+�����ӊ3r�p7h��|�t,#8�5묤�о��=m��G�؎H���g}�VXYyjL?��͛�����6��R���UcTO0�H�x�ˊ(��\�s�G��o�`�<���������`�`�5�e��,[0˾{�)��3���]c���/��s�J���(&�뫾{��BƮ>֬�
���+~Y��`:ޝE��+`�8&)�
�޷� w^�J��)kl� F`]N�;�l!`uU��󚺮[
Xݥ%��u�r�2�)�sK:�bkC��i���g����%�~!����7��7���5 �j��m�����;��b�GP���փ���_���er��t�	k�<��K6aҫϣ���O��T�H�w�s�� �)z�oq�ߓ���f��2  �c�`W��n Z�ԫ+���&M�' ���,�g1p�^�6KS�؃eѦVo&�6E��PR��[YeDǠ�p��#
�;D5����q�6g�B{�'\wRΨ<U]�P�V��q %/��>� X�*X�%�XG��*����ML(��>֠��jJ������u����+>��m|��WɄ��XO9�D���:m�4�D'��
NUv��p��=C�ҥ�镚O����1'[V��G��������n��G��cS}Q��t��I���.��Z�,5�N�z����q���pW�Ӗ���q	\[E9��H&2P�l����;eܾv��ه���<��M�YSŘ8����F���N8�Y_{x�\��/�a~M�Q�jR�a�/`�����8����<c��8�2V�2V�TzZr%)��KT���U��m���#�U�]}�
�\���Tp|�(2R�$�Q��f$�{:���\��&t��%������ƨ&�L&#�kB�� ���_R��s��������Ċ�g������qHo�Dl�4y��b��#;�^*�^#�QZ~�-�m���hO�2��Y�f�z\��T;GM�z����9L �ӄ_V��;/���c�} �B�)��3u^����`���D���C��,�"#`Y�����1:�"���go빨�U��h!�|�X�*cM'�V`
q�٧�Wvη��r<H�5�������}?�~�R4�v:AX��̖�ڴ�/Qc��6�Y����m�ĉ.��L�)?	���Fؤ�`4=Y�h�y���&��PR�4������OlQ`=��oۮ��'���>�@%�J����R�ۃ㈢�)S޶g�~��UQ�V���4����(wr(��5�0����OÁ3�oR䔅�G7G�&7�����L��B�F���t4�f��D�Q�E���%����\e�M$aB��!�U�[KM���Wb�z�9�}�L[���i�{�O�[�ֶ���*>Z�n�y�_m�E�a�Ч��P�7|v32x�Xo��3�(�����[0�k�VW.'
�^�D��?�OqKh���k�ѼC��j�+^J���,B�h�S�y��)O��
��@M4v���]�ҌTp�]��hļ��&x� |	����o����ӑa��<������{�A�v��ێ�{���n40h�f1���;a�N�	���4۝<b/�����4�����.p�����/�\�	��mJD3�t4$mb�dA}�ݔ�:
�q��	�>o"'���%��+{h6�����sB�6���)�ǎ�=�f��\��wf��k�Z�|^X���7 ��4��MV�'ňH�}�㪂�^�h�{�l�XՋ,e�{O$h�\ʞS��n#:W���!w֮k ��vP�Ņ-pPV����s�>��ѧmB�? X�����#>��/�I����ƚ[��4kP6R�<K�!�⁶��_���;`Ќ�@X��frR]ל>�wE���p+�u��P3��-Zl���s��j�5�A�8(!]ly�*�S���c�J���DTre̟�x�@��^_e��<��<�5TYpx�}U����7�=O�����DT�y�:�\�����;�d��o���P�x5{�8�j�U� ����27��+c�(�O�@K�����y�����+��K���D`�t�@U�`պ���vm�b���nq�TB��31�;S�Z6|7�P_������El��߳]�ANe�R3L���8K��;,���M5��i�k�X��II�=���%�Կ3�    IDAT]�����7 8w<��=��T�&)�U��nT��Iʄ>d�r"�R�����N���)�?2�k{��
f�My{��g��3�wz\.�E�:/j��g�6V�"V��c��:����<ƭ���.��Գ ����@9����:|�ґ�F�� X��� �/�Zk3��'7�f ��'f�5���)�`i�nE5�/:�z��/r��A��U�[�"��9J0
�K��ka]�أ�w��n�"��x��������M���^O�"�L��b�a՗8i8����{#/ ���]r�c��_6W#�x��.��O��2�X�;b����o��S��m�Θ�*0�i��1����z�,�Lћ�?��rYtM}��������\ �I�,x򧟇��q��l�0�z�X��� ���]px*�^e�%����+���7�����ˉt-N-B��(�⼴�~p�wp^�A�] +�&.~:S���W~H�r�:�dKlϯ~��-
�,h����^� ��!>�q��kd�o-&e�"��"��;�{����#�������TDĺ��f|��̸�Nd��,:[��e��T���%^*:��X�
V��KU�
[�kW|m���~�eK)��#`�ηN�����A��������"���L��5���l�]�~l�tkì���>J2���}�*'}�p�����P/ �'M�u�k�yfA_�A�6�� �4�Rխ/��L�x�PS6� �|ͬ ���W�I5J���:�E=O¨YI��X{~���!3���M�I����5@*���~ZOIO)?�D�jϑ�U�<ת��e�C����Ͷ�wA�P�ӹq���iTp,a	/D�J�m�Z?�ظ��XUc����Gd����MXݐ16U��U鼼�S�5]���A�1f�}�
NRk���8x�+�QK��>,�]>�����A4-i�M�^�͓;F{
�$��B0f"��-��^c���(k�B.t]�V"���媢�J� �\���e�*B3�P���~5\���&ܠ2���׻����VTv��������Co�E�^�v`���X�f�zt�t�]NkS��YX{3���˿ke(�X�s1��Ġ�6�˱��
����)x�;����K<5؉�B��ⵌ�i|n=X	XU�� ��qm�ϣ�<���mܸq.x�{M|�q�F���kl�Y�D��"t��n�)'���92 ���(�R"AC���v��ߴm��Ow,���BԮ8��Xt�S*Z	���Y{�u�b��x���&Fzn���,��<m�����Pc�ظU>6�Ӏ)e�X��S�Tybc+j]dwW��3 ��0��^�˴��i���chEĩG�#�~���Pç�4	,�զL��2�8.Χ�i���K`����d=�)�����V"e������pc}�z^��\w>8ۖ��K�X��*�ɻ���������tB�ꕌ��b�Gܐu��{�b���,_�P^6iT��@��+���x��U���G����6:ȗ��F�2^�֊�Q����ǣPHCW�kj�޳Tٱ��EwȦL��Ȳ����W��WM�Ho���#��ac�A�6�9��x��!�|�������������?%��HK��ٙ�����o9 �To�����yֿO�Xgb�����c��D���V��#��R��~��ޕ�����b���@�#0�֔��=��<��*{�X[���ӱ���d�q(c�	���FBqL�gL��>�7�&�X%^�d(���ˌ��3���s��ܠ=��͑�E�;Vy;�k��q��<�l�~�tYj�I��JY/P�HP��kP����D���Lka����KC��?q߿����	X�&����<cm��n'�w�΁U٫��v}�O�2E��<��z�_`i�ū�v}O{��h3�ҟ��,�6jjt���!���Iw�R� ��Q]\~��n��Kh�	Z$4]����H�J��,��O�kx+c-*�5��5�}hCkx�pL����O�z�9�j0����|��6ml\]G���Ǟ��U��7��n���S�u�ۈ���o�����R�u^��hȞ�M��s8��$8����U��+�o����Pc�dOo���nN�(�6y��NH�����Z%%\�0<���Ic�(2j DQ�'q�@����T+Q��ގ!I?��RrK�uPc=�#�!��v�۱�*��o,�����^��>m��?��5��ۜ
F�t����b2EQ��E֋/��3�vj�����&��Q��c�E&��GwP�s�5��O!���01��B�u螽��JL���5�,oh���n�z_e�C��U�k��q��FKCk]:����_��l�ߊ_�l�p���	X;j+m�6����]��gp5��D�*�)���H���Xٚm�=��ۛ31�ü&��"�Rtcs��"`�A��;�B�9뙪j�X� :U#�A���	�����=�]��!go&�Q��O��J,�s�s'IT���~��P��WצE�7hhԞ���d�X��ↀU�K��}�8�m���n��G{2�nCc�\�
x;�L�*&P���s���{or��K�&^���>�j�u���<�56�`�	��g��}�3f�p��L�u��q��d��E'U�r�^��}'c�:<�J1��D���"yN����Y�\p��S�˗�LK��DxC��U�V��L#��zm��4��t\>���h��Yb�U� �Y`I�{J�Uu�<" k����{�՗�C�9�ߏk��S��ݽi����w��hf�������[3=>TD,3��ë V8��5�s��e�}� ��g��Z��W^��5�MB�D=k�u��N;�W	�`�"V֪���>Ѐ���_C`�Ρb������$7I��Sk���3ǡz]�2��;̯� ��W_v��R�X3z�pU���Uvw_R��s������[��+,H0�A�ΘC|���lD_6j�Ps��+1�ӗ������+K��Vv���{t��^Pޥ�LF�V�Xc�55c���W�����x*��Z�%&J�]�����S�0_�%�o�$��PA)�e#
չu=�M�0���ƺ�S�z}�E�r�`@���mD�(�h�n��^�`�K����� ^��w/q��ɓ_�ŋ�������c��%�[��
J?�	�">�xi������N{~��
Xw�'�A��K��zk��R<�;3f3�������l(�bEB��o���>�=?�2��r`M�ΰ��M�O�\�QgI�.s|�)��kи�S���Zq�xܤ�Zl3J�<.|GV�x���3���҈P�(���+ӕP��D���0��fA�W��,^�[�|�N9v[�Q=��z��u*���q�͹6���W]p��]����t"�G��IQ��\p٬e�T!^�Ԗ�Za�C�/���w8N��ޟ��S�:�4��=q��t�H	}��c֩���I��5'P�١O�H~7f����|�q�����k*��Lyswf��S�!��������.�k�]W2�/�©�zW��6�{���O�e\���Ɣ	Zs�m�y���g����]1�9lԡ��c,���B�H�0� wy}�=��[�<k3s�f��"5l��L���\��%^�N{_� N���0cY|/��Tz��ZͫU�vF%'$7R݋��((�s`r�.�(��{��)os���in�w
���>
�ԏJ�F�fMC�520���@Ns��>���!0��G� QZ�`�b7��y�N�<~�x?�TKð�EZ��s+�2h8<��v������nRkkM����	�񛜱z�8� �u�G�n�;��r��g������-�.�zKvV�{Ĉx ҩ��g�0[�6`���UbK��V����:� 3�N�d�P���5ɦ�Ff�D5�u� �{�{�H�������L?��Q�@Z��
.9���0�9Dz �Ѣ�\L�U�z�٧ٸ���=w?nw�q�}����Fؽ��t{�eT�,�s�9��<��4e���nw�61 ��lj��-RX�3�u<�J�g#�y\d�|N����^~�MS	X=
��R��1�K#��֨�����Z7������m��X�K
�I�t�xI'ô�S쁇f��;���с��s���K��-u%���q�$;"+�+fG��>��V��f���=G'��u��?�-�S�7l"خ�ȵ��c�<������5Js��Kh?	}�ڌðo��Ht����Tc�8�򹴷��(�UwC!�z+��:0q��yt�%j�$��Y0~�&(����Q�i{��z�C�!6�9��4_[c-y��L�HC��|�Ջ���U���m+�of��� K��}x������sG�G��q�)8(mks��i$��ܞ�K;�8�Jʊ=�>k�k֨{{F��6=�L����:�FXc��z�ɧؘ1cܿ�����F�mTv��~��6�؀��ic��E̱��t`¿�d��v�*A�ql���z�׏8���;���,{d���?8m �jiN[�0�%�v�:������/�z��^�4VZA)=N �;x��F3����C-ō�`�JX7R�8x��j4��w�y�0��և�IO�ؽ���=��L������[��C���/8ɞ}{�]��Zmf1ub�1IZ΍-`�
`]�������_h}+��*x6S�
�J�$*�'`��I�����KZl"���m�����#xF���6��QQ:���l�1�T�j�GqDg�AT�C�3�FZ#���t��Ȅ?d'_��7�lͿ+F�I�Xɔ'�ڸ_5��v�";`�]��c��O�W�Ks�^h�:�0��m�V�ڟ�`� ���>t*���oե8�:Èf`u%��_���r�weG~(�ò�����B��@�y/�L4j�''>m������ocB�ο<��9�2�?�S\�t�s�%(����k!���t
Z{�ч�x�{���lM��[��U�]�'�I|����N�^k� ����ʫ�k��6�<�x w��=k��52�]��O/7៊��1�<�w;��M��٭�>y�����u��m��E�������N�����>@|$�cY�7Y�=���g�P��8���و���d�ǜn��Z#>t�������]r�4.���ƿ�{!v�T����'�׮���n�΅߶���f���]6���kuDߥ��R;�$!��V�|$�����d�좁[֮�o�kW�} �H�GUг�o��k���f�D{�qٙ��WF��O�k7�'�*�@��R�k��T�-�:A{�;U��_�[A�"[1�mIjl@�
��y@s0<��Z�/��DQ���dST�[���ӱŬ:*�e�x�q�ypk��?��T�V�BZkA��ǚ���K�ROg���S'�8��{�ik�
��(��Zu�,b\�Ğ#鄋g�{o�~YM���Ւ��\å�X�F:ORl��gVe��}��@�&`�e?����S�.���R��^bc���|��v߃��B��� ��@��Bor��O�7�\lw�}��˪|z�%۰(��g��QTc�d��4���dSoaO�c;��Cm�����b[������m\�l�u���FB������ ��W�4j�i͕N_��/��3g�W��ݧ�tQ�ᚊ��x�v�y�ꁝ�>��<��!;بC��� �Yg���%���gw�I)uٸB��Glkx;fs�gO{��h�Mq?ۓ(!��6VGԐ�ɬZ�����ևz�.��Rl������\�>���g;��Zl���j��U�[i�6����?ؼ�k�
<Ap*���+*��o5�w��Vq@}MDMt�R(_�����i%R��,d����L��۩���?f찌��ڋS/���Kܥ������J2��l)x��P��� $��	���7ŁU}�]r�g�j��>u��XȚqS2��m3�z���j����w��e���A�\T��g�#v��U}��n�e��Ͼz>�TPճ��fx��%�	���#��Ǹ�a����zG�*7�,J4�b��������8��]@����]�#��ϻT'�J��D��-*5�������l�@�)�;�P����ٿ���1o��ӓĨ��^�����]p����}�챉O�i���~���p��l���P��K�\�ԉ']�(���ٶR�-��H�ܗ����m����&����v�L���,Ye����g�V2�r���aC��-�w��v�=Q���J ���;vR�����Q�m�i�6P�[<c=�0�FT�xmy����nԿS��������*�u�;o��J�k{�]:ڲ�o��/ �~�A��?9�&=;�nA uՕ߳�w�������{+�o��Z��Ŷ��]t�iV�$����g�o;Z��������[��|�z��9�}��	
_���7��vM��V���y�ޣwd�#4ϩ���I�G8.�~�c;h�}�OV��]��^�1�Z��Ҏ#���E=�#��&���B�z+��,���d}ț
X�k0��`5�Z�j96f���XdD�˖,�B^��2Vw�ل>֞�����V��It�T�C��\[-Zh�L��ƀ��@�K���
��җ���^�-qd��K�)����#��պ5�m�Ww���D��!d`*������5��aɺF����t��Ͻ+��2Z܄y���/�)._��qm� bc��Y62��`�'D�?g`��Q����v������wf}� 4��.50�`�j?�Gv�q��l��Գ/ڣ�=�=�ju��^6L����ʩ/7��?b�����!\���}*֯��>x���LOjtx�4`���_f��-������:{��ќA{�IUp*�r��*cm�,9k���4�5����/�6[�
>��}й"~���{/��v�3WE	Æoc��X���E�UY��k��r�V:bg��� �Zg�z����v�o�|�v�N�?��=���v����^�m`��v����w��w�fM5����ng�}�]���2cq��f,>eQ5��9�$�h���%��
��r)j�W��B?�^EŊ��xR	gZZ�V�74i!�Pu;J�����J����*���.^������� �&tz�r��E�]0�LژȮ��)T8�\�b�X}�kt^��fKl^_�k��O����%)�nT��(!��m�QH�
�,�&�>G��A�_�����w�8��)3Al��4��=wic����[��%+T�d�c��j�����xm�=�س؟b����I�j�}[�����\`u[W�@�ns�,�p�X�8d;��C췿��ޜ9���t0Ȅ�ltqc�JX�j����=F���&/�k~}s�Gڨ]F� �bA�ܣQ���2g;����7ޱ�f�ğ�VH����W3��~�o��g��_c��T;epm�+��\�N*x�=��jl�9�>�;M��}���@�2y'��I���f���F���籊
vU0�6�J�C�U5V:_�h��ti<�1_���@�k����+2l��0��}�dzM|i��E��u��f'[�r�U ���Ϯ�������,�����E�K��D��.��v�g�'}��!C�������^}�#{m�<{}��)�R�=���P���IS�l����"Y�f�jQ��US4U�����*�"���E-�h��WD��Є��I?�%i�UW��rm�4�*����|"ż�m��X."3�0sD -��RX��f��dlJ��ְl�1DU��d�*;h-�������yI5V9/��J�Z=��/�K�s����V���Or����>mc}H�Ӈ���Wv�>��{U��4$]��&��U�(רm$���
�M=1⏠�NL��d���L�7?c�ЌS(�f2Q�#�P�KK��1���3�8�~������/��x�#��ֲϮ�}�e��|�`�"tl܀�e]u����$96p�@:3��P�ש�1'�9�&M���в	��#N��;�1�����3Ú=��5�ß V�}���Xq^Bi�֨
����=[�ӆ ���n���*e�^I�������#�nx���K�Xc���X˖-s��Yk�QW<�S��H�"�%q�    IDAT%�z!�3"h������1'Y~���t�*;�֊�O;�^{�#"K6J.��|�p���t��v�Ï�qǟA�ζA�@3wNf����>dh���a�=��,{楷 U�Ґ�Tm����*�d�~V��Zo�][=7d��(L��d� Cu5K�Cی4\�PnJ�1������B9Y���QXQ9MP�d��nV��0 k����s4���5?��!2\Yx��DT���+c�P �X5q�;����DU��<�h�ࢃ�ހ<^���;[F� o���/"�~`�RGؙ�&��
��4�
��2��f�E_�	�����r�w��*M53z��.�~�-�U'�Ha�iѠR�z&۹io�O�鯳9��#���ڡ�Z)Vq��bn�l��
>����[��gΣ�� ո�4[�d���s�]~������>`?��O�7�5��#��*z�6��-,p<�?ɠ�Q̓t.��V��GW},�g?�寠�	�l�ɞ2Q����ս�k���
N�X5�F�%:�,���v�l�X�>V�X弔K���#N�Q�$`����S�}�	R�����:(Մ_nc�`����k/���d�Z��_pl���H=���c1�֬Zmsg�c��	{}���T�+��;�z�J���k~Se@sc�p�|�K��W�]w����k��h�P��f��b;���섓�����Z�����zsZVǓO�N��l2�V�
Pfe�,�D.,��4���"鷦`�\E�]��h�[��"���nX����D���51,HǠB�����>DZ|˝�X�4l���g���Z���2���"Lӱ�@�����C�D}��F����Q�{�]7��kl\l��"[)������F�Z�Ns���m�7/�p����vّ���d����i�$��Y(Zu��&6�C� �n�� �^��l��Ȳ<���з����&)�z��zl���4U����ϧ	6���u A@���/��SO=���{���V�wo���j�~p��ܳm��v���S���J��?���b����=��UV �+ё���ƭ�'js�JIl�iR�ĥ��x�ܮ��O�|:t0�H������%T�B2��=c�*��K/�vQ��?��{*�Z��j��^��iй�*zj5輎�6yL��e�I_��+x�=��O�MP-^�l��=�Q��<s�Gt
c��~�)[I��z��:��iC�u����S��;n�ޜ:�e�d��;�;x���Cq�y�&��:N������*���C�s�M��⥕P��\,@IJ_f6Jq�Q���	SU�>H��W��ںLi�^����jcHф­P�t|^�H��A������,\74�>�&n�F���`��Z��λ-��āUk=?V���s��w�&uك�8���Y��2VY���S`_���{�hN�7�z�C����GC%�ڌ�KY�j�%��w~نwn���RsfA�k�(%6���>�F^�s�DM�֚ɵ�5�t�&�wS7k��)���t�^���G����������0%~7��6�	�>��7�5���c��iIڹ���x�t����dโb��tߪ�D{�ܙd}��#�z�2V�R�ʣϴ5 �j��M�=��t����od��X%Tr&Q9{��W������X�O�
���mV[����K���3�qҍ7��m-��V�c��.;ۅ�n��1����c��̰���~���ދ�?���[��љp>�h�����`���5O"M��6�YFb"�c��Ŀz��P��i>��*:W"Z���λ;/��u��l�;�<�U�*��\�uS3�~���L���7�����oYQ2֘�k��bK2u����z{��'�����D[�k_����*����Tu��֢�.<�bb�,՝�ي��ƫ�jukۓ�q��Õ���<[BTԬs\ 1o#���]���w��"�j��z�P��iv��p )))�����i�2S�k&�kn����YL�o���િ��/��X�.Q�Uk_�{w;��}���_����sQKh�	�\�;Ԓ-��^v�7O�gߘnϼ�:��мrQc3����
��8�`�����i�۴#^R>.*��#�VSW��T~���D_k��u.dn�=a� ���x�S�:7���0�;�a�{k��ˆ~7��L�P�J���ƪ4����*����ک��J�t��O��������WMP�O�PN7Z�
�D}e�qf�d)�Ų�j�
�`u�x�<
\��w^G���gb|�5^3h\#�ƾn�ܧ?	��D��d�z���׍���2�("q�K@�;0��%����t��F��#�P���p^\��U6t�ی�5ڗ�3���|��2Jp���F���4FZY� HI��{����uA�0G`���JN��al\����7Y3I@.JV�5i���HykV��0b��@���i}�&�aJP�޽����V�X�^��\���i`����m+Ak�!�/$�`QmKaЉV��m;-��aD.b�z���`AU-�I��w�Y4�[��\�<�߮fl�P��K]���5𵖌�ې	�/��9�_4��y��7��I�ӪY�5b�2�֚־�m�<��W����Շ��y ����ڹSX����zt�1��s8��X�H�|#̠�u���ۨ���h�%��j4`j�[�l�X@�\���Ҽ�Am�P��"�s����t9a�8��=l��ǈW�+�vXi
w����>H���"�݈AE��<�x;�{���+�%��&}b�nZ�)�F�}v���쳓=��v�c�h�E���_c���h
��݁�C�us_Ei�=���.X ҹ�y�C�E��f�Qu�Z
�F���2���s��0}��?�����iST ���$��0���G!^nk[X[�'m�[7�*0��A%�ٲ��4��O�l��|s��d�)��p7��S�6}tt ,����@���פ�D� T�u�f�!�u�M~������i�	����OM~]o��J�=<7@ox^ Ş��5V��_�|>��AP�SP��X%k��=f��d7%�!�v�J3f�+V���
\�0��ho���J`5�Տ052��l�e��_bs�U��*��]/��< ����d�IT�`���=�}��Tm��(~5�5��I��5�Ҋ��c��1slT]����.��o�d�9P��nto˸���3sp��8P]��M%[��(`�X'�����\�o(c<=P�uY�\���ںY?$��
6��f1�c��O�
�h�i���w�Ɲ���5����u��n����5;����.�OݤS���J~�R�′���Ӝ�	�Fq��QF�nχ�  v�_~�G,�&��Ū��~��T��-d�����,F�>��D_R"��3�'�wmd>�5��Ye+C�;���i�<�N?a?�9�V}_\3I��zV��QE e��'�������� �~<�.�^Nƺ��q �\���1c�^�Ё՚1��r9qX7�>��i������ڒ��zww2jI��5�7˖�b�i;K��W�-�#����"�N��K/�˯��5V𢡊5�Zz%7�Da���V`ua����`i	�
�-+8�,��tN�s��"άxX�B�vf�����jI�׷�Fg^��X���g�X#�P��U^; jؠ�#*$mk�7;�Ք�
��Fqw��;�-��8�:n�N9|�����8?ێ<�p;h�^��Ģ��Tk�3-[�~XeO=�����A&�3����&���x��rܑ��Bg�n6����TG���Q�<�t8����6�MB톲�4�I��@�]�ǃ�����z�n�
�%�����^y}ײ��YMI|�٣3a���V"e�M:��>�us�(+f(�+�4�C��
V�ए��b/����� ȇ
�$����l>�:�E���y�o��O��D ����I`^sLRGk��F�)�U�'c��� �<;�:��q�PV�G�E�F#���q���z�p.��w�|��ͤ¸�C[�$NT�!ڔ�ΙІ�
+���"k���O��GV~��k�Ԯ��:��>e�$��UԔs0��2��fm�C���ϰ�4���Y������> �ԅX�56`]&*؁�܁���KTp��V��t��[i_~����0�,��7�q�`0 VQ[���Tk*�8�g�݁7e�٢��#`�$�`M�]'`}Z���t��UK��j�C��� BK2ly+����9�+:����`��;�@�77�d&٧@��5�mɝô��v�Tj4�B�f�a�	�xj�kU�X���`Q�8[5 ;٥��Ft*랍�����X}S��5l�]�ߕ1wwB���v� �I��w�9� C��F�.7�駝d�}m����,{��W�"U�����	x�yE��?>jo�3�Jը��5����w_�	ͼ�cۢ7��^l��5��2Q�������IQ�>�Z"���C�� U��9��)����+X W��a����;�=J����c��os&��`+�����`-+`�釀�4�)���qz�t�Dgi�_ʊy�9cu��r�b���f�ȁ
���S�q��1�jVQ�5P�y ����i�Μ9�O��5u�u�8��_��C�+5�f����au*X�u�z�I80����l��YrrCۄ0��+1'9���EISk�	��(ϋ���G䡯J%�!�&#:V�f�R�o�b=ad<�ƪG$\�L��Y@���������'�"�{�}V�D�@U"\uD}��C�o�t�=��"����O�3�.�ɦs�W;�.]��=�Tp*��[8́�WY�]xɥ��<֙3f����P�d��~߂���H7TOMe#��at�T���p'KC��u#`���[^a/W+c��%~]O('E8G[%�
ؒ�J\�X����SX�*XCM1d�->-$�n��g�݊���t�WWV�w��$c���d?u\T��/]]��>�r�"��?	�:V}�.�V����}��f���<��GJ��������1�|��>� ���L{���C2�0��@-��_^�}z����@�������V2�G`�����T(��/��u�j�!��*���I��Y�a�U ��H���rP�~�}_m�q؆�W�������a���K �������xH�x���DT!�J9�B��-���1�����IT0�6Y�հz��#��׹�b4D����j��ޞ&�s��]�t�9)���|�����s6Rc=��=��1cl�xIّӺ k*\?�:?��smԨQ��[o��z��Nt*Ō#k�خ�����L"��3���u�Y�Pq�e��֚���%q��Qe�\Q��rN��%���&��,�L=p�QC?��+��>rZҬ�Vd��d��,5���X��qjX�@��L��4�|[
��m;��#��>e4�/6O�H$��]F��w��ޙ���,Z��j7�MJZ?���`��1�Gl�i(��|@��N`����0\�9���Y����5qGf��抗Rk����!F��У{6o�T*�!dJ� E��V���O�<y�����:��p�N��֥kԕ��3o���3 D�Vۥ��4��DkP��j�z�x��j�DBWOXIt�M��<O�v~It� �������:�xQ��Xi�<Ϥ�[�i�xL��j��j��m���wu�8#���׵����R�> �������8&�|���_��}�E�0�ќQ�Fج���o�c{u���׷ѭ F*�7��/$ r��.L��/鼅:�2U}.���ϦF���I�>̩P��6��ku������1�}_�ˍxT�Kyt��/
��J�Z�#]̞(+X%$!c�8�.^���������U�o�s��bN!KC���/!=��L%�}�u�8Q.g�<��:{�<$?t�lbƚ�1�Ҫ���3���#V�4��I����'�|������y�(k�F�A�Yl4Uw
�O�e徙/�7�VU3��q��C�Y���>"*���9\�>8dW�Z�\=Tׄ}�F�V��hC��m`[e�`E�&�|�q]SUcKqw�w�L$T���:�p� �q��߸ҡ��zԄz�7�&�i�8�������@}�t�x��֦ZNY?2jE��}����J��M���1�j��4���K��.���- ��fџ�	:�K:���Rko�#���]������x}�vSo�q�ߍ ���r���q����s�US@w��p�R}F���X#��ukV�~�7x�n8D9��3xXUk��c-L��dw!;�_��Ekp�LѨvO�:�(�x�"U�Jd������:��UF��1�/�2TML?�⩍�?�[���6wm��.j9̂b�3;���U�:��X[c_?�H;������r�}D���~}���̇S�޴�9�o_�g���knǜf��0STiL�qx�-�m�}��T��'P�T�2��g��x~��5��^E�M"Q�.=@�bY��'p V�!�GS�f�D�qmw��p�~G���&8^�
�r�$@M$sҦx��~'`�`���Y�Wh�'���o��Ꮾ��Y�|�u{���كx)&�X�����ޟ�B7,1�ߔ�6V�K�n��F�z������61c�X��� �T�����sζ��έ���z��}�M͊�I��Mr���]̟7���d�9}Pb�jyw�5H�E��k�v-�z;��v���fv˟�۴�˭������U�N�*�b̘��s�e�������_��&Nz��P�B%d�bAu����Z !�����v�Q&�m �{���n�	�����	��Jc�x��\��h��gd�=7�}Q�a��g������K��M���$��n�z�ŗX�{ ��g���XU�TX�V�yn��q�i�ц�?�[�5�H��p�v
��w�I}���Uǧ�uذav�a���&�|���c~��K��;a1�"c���B*��p>�2;�e�KJ�K�+8j
kV��?N_zE��ЂԦ��l��&}B�NN��&gy;���dς����?�"���z���{�&]5�l�7�d��k#B`2�.p�C�Е���N`����~̞Cp!�B�Zm�lW]q�؇Lb���(e�*%44P������W>��a��O��{x�}D���#3�~�P�N�f� KK�Ϩ�)�	[Y�zۍ����w8��÷�;3��k���Q������Y�b-�=��RWE���U!�X)�EŊ�lð"K�L_k`\t(VI���Y�ڿ��,�����ADoz��:�4w^Ҡ���ǻ	�ʌ��>%cmӸQ�b\���C2��ظϒ���m����X=��, ����c�U���O?=L�Y�`��H)cMU'��z_b�A�����&���Y���x �Υ
�0U&�K{c�:�?�~x����f�ɛa3�|h�1`<�]e�m���v@�����/�b ��V��D�hl�Fux�.^���6zUfF8�8�&�l��O2Ɉ��T�Yf�w��{�?��t٤
����մU������U��\GdMH4��Zi߽�"[Ɉ�?�v�S�rB�t"���\�!}1�>���]�$*x�����^p�MU�N�0��8�]�� T�	��U�~�Ծ�x!�����ͨ�I���l.��=bv�����:fm�o��S��L�*X���W�X!��M�u뤂C���&zmn~4�XkI���y��iڼ2�ٓ4;='[�>��@�6����O5��� V�2T֟��4�Du5i����9��j��P�37��M	d�k#�� ���
S��s�\������t���L|�$m�k�RǦ��>���Ӧ�G�>uϖtL���S�5%c�y��X�2�o��@�Y�g�?n��f΢W�L�K�Uvv��>^�h��v�-YA9�m�Ɣ�2�����uk�7��_�����a�]yť��hk%6��������9\o~OTN�>��q���Lgl^;נ���>do_��#���C-+�����t�͚=�σ�M=�+kl���LSj/���s�=����l�LGL�Z����;x�5˝�{λ���oC9�����E�{D��]�$u+ػ���^����9>6��f�ظjh��}�*8�汖�*e��n��c�rZ�ʳ'<s�di�e���3N��|�+n�.�!�{    IDAT�c�c���]���fk
X�X��5ki�)d��u��w X�)�W��Z��<� ;����W���9`��s�W���k�-DT@cq�gF*����b���'mnNY�'�Y�P�շ��|㽡��|�b��R�T���[Mr�gV.J�6�nX?�y�� )Yi=�+�+�R!2*���c;�8�7DU|�=��.ԪD^��@ҭ�ČÂ�z2V9/U�n���A]���D`ͩ}������*��.���m�Ǫ���ɯA�� ݥB{6�e==R�O#Py]�{��C٠�x�6E~�xݢ��o(ʂT��B��Q��!��&�f7�G�3c߀�裏��&*��W_�/5e�A��X�
�����n�  k��(Jn�Y���ɡ��N�eB�9'�J��v~�kK��+���kk��Z�zE�����gr�2�Lҿ�͖�m�� ���L��W2�D��'���{�~pv8���/ (žn6w4�,&�Z���6�U�oH��?U�$����A[7�>��=�XCm9d�z�����597!�O8 �k���#	�k+��n������׶A!,QHb�ի���Ys����D���[��oe�L�»���(�u�T
�t7n�'kVDd@�� B�">XE��9N�݆�-��\v�ь`Sf,t��� �U�aӦ·zĪ<՞O>��� ��	6����T}�k{�N?�({q�<�G�<���<�>�E���~_�K�v���.8�봋?Z�=�n7�>�x���w�_lM
�,uQjt��������\h�N�t��V^ޫs�l�^�ZSC��Sg��I_A���wr~���ƚ�xiS,X3�{��	X=������N�U����3�k8p�9�>e��>�����z����6�*D�uUDS����]�N���ڮ�v����*������������wD����??�ٮfK����'���~�Md��Z~�6Eբ��L|��h7���m��,�Mć�r���V�Y	�T�a%����6�?h�~�h�4"��{�շ��'^fض"<
�K���k���K.��V�W�S�Iw#F���ݦzѻ�e܇��]x��X��*�j��E3m�z�QS�5��T5�,���g	��YQb�!f�����H`��UNW������x{>�?#��諎QT����`��u�ԩ6��{طΐ[��$�z���5ԥ��L!S�FآX6�E�"����k���r�JZ����<���F�Q������U(t�դQ�������k����#�l�%�-��i]��SMD"��H����R�n�� 2e�yh:��c� 
�;�aB�*�@!lh�A]8n���_�Q�=�4腺p2�B���.`��c��W�f#E�.<���=��U�H�ݝ�V�(�tW��ؒ�?rOn�%l��4>����8�����@Aﳵ��R�Uk[��M��+ί��
<��ϕ�¹�0�W�_b��|�3���G����G����.خ��|�n�>v��w��^�a,?��%�����,Fg�ɌGٱh]@h-h5!*;��g���__s��yo.{a66�c�t��?������;�_֛{����/�z��Ly�F�F������6��* �jk�X7XU��nkh�Ȭ�t�VQ�_���:�u����!S7b��45��+��6���g��YYf+��i�(��(��S��?�m�L~	j7���m�G�5�݄�B5/�����]vE��0�����Hз�n��A{��t��\�P=�"�d��٬Ӈ��sP��A�M����a��É��6��1�˶<p�1��gNx��1����
kc�y���H�Eݙ���(x��������`.�b�G�^���J,`�xI��{��|,�W�emP� Y�څ�eקWj0�YWKο�O�����R�-R��+�戵WѾ�N���ܲ�2�\���f��\�{��~r~���Y�2�~��g�{��5q^���֭���χ�_A'WRuT9,��j�d��IH.k"s5�\c�������ᑥ4h��t@}feY@s*X�0	�U��ea���,��]a�L��F-K��Z�-r���~��>ipb�W��� �مJ�mD��Bk��Xe�!��:�՞�F���P*v��8�Z�Y���q�Z��~Z�DC��K#��ztp�{�S���6e2����5(�5h�,���7c�2��p�{��l��X5�Qf���b�:��I���I{��!E--��A�!`���X��Q�������캟^j��N���t3COJ�o�r���ow�=����kVRZnm�d���vх���k��3�N;�wE��&����C�f0HE�z3�Ű���$�,-ʳ��wm���k~͜־�����kl��vݍ�X>3`����l�s��vf��16�z}*��d�Z�qй�`���*`�*X���Q��/�q���t���:3V���v���X5�F5V��7���n��<p`�驱�(��Pc���ށ5 i�vz��o�M{�&���s*���β{������H��{ϩ2-�z֓�Rx�ʷ��Ol-~�?��-��7>'T�7Pg~"�8��([�*$�&AV�[�n����^�ٸ1{�V3O�Ui��+S��g����|�����v��E05C����G����y��x7�o�o���J\���.XsY���֐���[��5\-Q@/u�C6�ZQ��1�?�
��`�h��<��;���6d�T0���q���ާ���zG/�Xo�<�G���	������r�`	QV24^�`ykl�T��4T�ukW�x��:� ��*м��D��j�@ՂRQ�J�p��z���P��P�YwŦD75��6�����>�Aa�7����*�Qf�`W����{mI����j�h���=��V[r�챛��)*-@��k�M��h>��ze�kO��~�5�z����F��xMQ���EU���B�(�����3S�-ɸ;�qȈR[n�ܐ��P�־��nvƉG��^�z͓sW��>��О6k�:���Z%��T�2��-FAba��Zj�
`�D�x��~6X}�$�A�����د�<�}0�G܊��QnG2����Ю0�@NdPJ+��Y�z�m3t��{6���Yf��_�eÆog}��-�P���u�
�T�U^R�^l/M�a�1	�x%B���?�ɏ�b���ndm�s��ܻ�)ւ�v2���'�`ĝj� ZU�5��X�kj���a=9/���n��y�Vъ���X�����X������u��V�5/�*�٦U�m�Q��O�>�^m.������QD��Q���^���W�y����Ғ� �8����%���O�j����b�����*�+��V�hp���
+�|��ع'��
�� �1�hm����G����#9EǵP�8u����0vJ�e�(��`�}(�D�����Vڻ��xeiX�����y)��UjK��v�V��O�ki�}�mԟ{�c�u������v�Z�L3S��������Z�׉ٯ$�
d���^[mT5E0�`�&�M��J&X��|ѢE�oMr�T�\'M�)���XWɵkk���`N�'���5���&�nQ�OG-��m㭬g
xn�hV֦��ڲP�Kh��C٢����ޞ�f�)c��#.��X"#�Y�j]��f���Zi�2>�L&�� fd��F��&lG���Uƚ�n���5'����iX���D�̱����k�ܐx|�6�6����<�BY%\Cl�ȴ�>iL��3�?X��!��./d9C��r��H��È!���<l�0Pm1p�E�>�h{�5؞}�c���w�Z�e&�ڐx���4�j�gt�'�v���?��ʳ��e�݁�j�htOn4c�5��ȩI�]����m��E�{�c{��m����m����t|�0�b=(�q��ë�R��W�ك>h'�|�1�f�[�D���4��=z��Ifm��{߻�&���=�ȣ +��5�:��.��2�x����X����D#��X��h�al\��N`:x�����M��n	`U��wv��op�ҧe�iL�A��=F�h�"6���y��>�U5V���DF:K�6���J���mU%��K�r����*���O���:��ђ
ۥ�}�rЍr�Ac삋�i��Y{���QG�ԙBhٷ�I�Mv��16v�Q�4�'&O��l,����Dƞ-�K|��)c��������":��#��'�a��O�&�+ ��w��������{�1���=*��\����D]p�9�����{6�z��5}�<�lF(0��J�v��r(��>�ɲ%KE���=�܃�X�gj�S7��� J��0���#���?�H���F�lU��j��.��E���6e�k%f�z)���>�\׌:`@��U�Z�[�XU�ٚ3��֥J��	V��<1R�:���߈�`'dz.�P�Nj� U;�A�m�PDKy�
��Q�l��Z���D eԯ����&c� �s��&%!�X)EU��iT-9(�[E��%�j�N�1�v���#֐�F���3M��JR~"��W�vrMSz��֢Y%�����5j��5�ںԪ	%��,V)���(_�/S�W<�{�T�����\p��r�J|��=�\�qd۞��f���~��LSYkoO�a������l�6XG ���~o����6e���X3hFV�������5���ϫ�y�+ʲk����R�ʇ�X�eǝ�W9sSo`�R&�4R���jHp�<����礧��3�:����ˀi���m��eB�_�{�Z!
��f������6g�*��R^���yyi���c>���~��\��%W�pK7�
��X�<���j2�D��>��mR�5��RU������c��rV{]{���'����`�Z_������v���4������
���ReӞ~,�t�I����&���xF�U�'C�z�I&5%���_ւ�]7�Ш�� +���~#�
��O�
������f�O<A���7>ԢB�W�k����m9v�7�|�s�v�A����lp.>�fu������o[+t^e�*b"&"�n
��8L&��bx�:��wp�R�v`�Si�ͧ�?�^Ր�k��éKzWg-������א�)���Y��׏a��O�����]NoV���lݢ����NP��(ʺ��A�,��}&-l#�8�O��d�Q��<e��/���F+J�D��~��YdSk�q���j����m��^�꧁��a�*����F��$ woj���]Hi�.����c�?�7g�qv��t(��o��{_��3ꇓ��ʐ����B([l�"���y�2��t�AC�iOh�/z֌7�U�����5�) �Ԫڠ�֪�>���,�X j��m�|]��v�a��<���z��y�t���O�D�!ɓh�b6W�ΘڔAOQ�"+�`l)�U��n���߯������W��|�ٳg�)*+a�P��o�!�������Vܠ��n�(�${�s�3��C����q�o'��L�1�P�Q�@E��1c�`cXH+����;Smڌ���~J����aH��.�r�
�"�k���7�����×k3�tT�(�j��)Z�p���6�!֋؈n�6���S�d�Xu�E��9��_�ʻ(ʰz<��l��"�������,V���_�y���v����lsfϲ�=��>�h��ާm�3��`Ѓx��R�{��>�0�R42���/~�k�2-�x ��uG��e��l�~�۞d�1�@$��=_�O�<�1T�ի����.��F�&*��;��l��c�ש�]�?���;�d�z/j�u>褩�{*x4eɶ|�p�gd);]�خ�����;��ɧ�����Wx��XXW4��m�J�Ӥ���k�������8e�#ָh5�V;㌳|й6:��V>F�=�C4���k�q0ro�n ������oY5M�V2����d�%$u��|��D&�^4W�F7�OZ �Q�_6�
�&��˙�Z��a��TK��y3<7��$7���G��w�N} ��S�I�\|m("Ҽ��A�ʚ��/|�Avֆ�C\�D!d��f��p��g��'`�`�e�e�FeT-���<��q9<�<-���
W3J�$0����ر�&�sWA�(`�Q_��<�(T��L:%'���:[�f���*�.�`��g�W�=oL��S�EǬr�����>1H�0�JW���ظ�LF��\�2��#j<?y�m�Y�|��j�&�h|��|������6WZI!�d��6x�0;��<��>����瞟d﾿ @(�n�&�}�ˆ�~uv/����4��k�ʐ���9�aԎv�ر^�	Liq	u�j�0a�9��:N���A� �+��K����%�Q� �5�\��V��;�#\��Ql>�����޳���mv�-n:���:5�U@�Y5}�ʹI,��	M ��[e�M�]�����B^=�1����倳�tr`5T�>l����`�=ww+S�k�_�%K�aL��d�v��k��1�b��Φ<I��:��Hv��)�l�j%�5����w����\�S(� �)3�� ��CG����f��>��dEѺ���-�vu�󈶇	�C��ϳ�s>�?�v;�#
����mĈb��g��)�رGa����u�3�w_e���q�Qv�ѣ������+^���ϐ潄���u���KO���׹�w>nvc���:{��/�Ӣ̃��a���u��6�﷣[Ym�h��袋��d��\�9���&u�oğ`�rZ,g1�|U6w�b��rc�Wz����Ïֺ��I�y��S<�P)�5L3H[az�c�^�����^XXWX�ا囑$�20��)@L��3�c��s���t.��ۣ�%�cA���DY�i��Jf%&����焽?w����I��!bؓ�q���!d@|�=�;�Ρ����t"��\Ԑ�N��4���ɣqm���S5B�� ���F��MWH΂{��BR�|��.�IL��i��U����"Ch����.�����V6͏�o�a�I���0��N�^_ޗy0�(�j�-�?݊8��g�{P�pAQI	�9:��/V6�0�
�<(���iS���6����Ӟ#��c�4�h�Z(�s��:�j�֨
��Wqk��6S��&2�j��HkI���9�Um,|6l]�.`�j���z��6{���)j�P`��И�|2�"2�l6��@cd�\�j�2.� ��p�i�Qsk"�^{�M{��<�e
S9״뺂����P��T�^3���[�t9�p��w#em���>t��σ��[S޲>���St�ْ!*�`�řc0G�B+BŬ�߆�S���aC�1���f	 Yv3���s/��|��o�+��֐]f��(�c��΢�lhV�fK�(}�3c���No��A������m�Q����fg�i��
�Jd��/�hU=-*�k��m�t�K���6��ܡ�Z��TT�O�N����a5n��㺨N��[�!�c� ��ȎB��j^�4	�u*uL��E�x�]|�>��=ؖ.]j��2ٽv���է�k�`I��ԩ�����]ƨ����������U���'N��u�n����W�^3)�e���z3uh/���n�3g��6c��kU"!'�����ҐZ��<�񻬽�cO8���tH{�=�a���;^��=�U���� u]<3��-cȶ���GZ��0�Q�k ����H �(H�,_Rۯ"���n�م�C����5���E`�ٛ�D����塲}��G�~�4j*�DFe^SS��?��.� ��+���6Ю���Y���z��kX EA��~��V��URcm�@g�ʜ�s�A_��U��yʔ߭
ۛ�üH�l�	�����s\��A6)zJl�"�"t�k�h����"�q1��u}�@:S�nr��x&�*b�����H�X������I�-��P-�"���������1T�ea{�� ��:�=�.���DeF�6^�X+��z��O��5�*�ɞM&�:�v��u������IkL7�g���q�(c�c�n����qb5�\s����tf����e��9gD
�    IDAT���� +h�1""kL�gp{3v_2�B���������-�$e�ȑ܃�D����ZfY[��7����)V�!���mv�mbU��ĽV}����O�;6l�� $f�؜�*� ����ΫZ`�*[$�*Ê>�{�!c�v:��t�4)���|������l�!�
�	`�G���m��
�l�<Ղu���=,տ�(��Q�ɣ�9w�<�.��,����J�u$��a�i�ϧ�Y�zW���� |,�C�1�#Ґ�w�@C{O������G�\�OR��m5|~]���JE|n���H.큀ց��)@���b�|}���+�y1���k_Pm]�p@�bŲ0-F��2��	�`�f����W��uN�{[.-���ٝ�=w�����]�^*fA�^��1����J�y&�}Q�� �qDL{�j}�XǍ;��5�N�Xr�	�й%-`b@����>ZdO??�*	L�z�}�8��a/[��nFy^Ho���	����Yj�K��*za��v����5i��z0���)��vo�����3����)c�����zj��u~É��C���$ʨ�N'77O}�F�ߋ4�z� �m+(��ǎ��#����{��P*�V�)p�@P�E 4ϻ���S6��p�E�&�&����ڑ&�h�MR
��,������C�ȝE&�x����f�`�v;Ȃ$q��~R�u�TY���w$�7Q��,:����<d�����3���� ���l�{����l�!���In �O�y��5��s�ɯ:u��d��I`-^%�{c�����J�(Q����-,Rmв�S�P�B`��W�r�����os�E����W�T��P�
k�_�)оm�H�AV��ռ�y��u�qZ�]X����-��M�t���*%�ʴC��[YEq�F���$Z^�����7�6%�{����WV�qRc��5������V� ��������޽{��+��}w�,�����U}K놀��a�e�>��� ������u��k�L��;)�,/�3�U�[{u�Bot�44���($ʢil�aH�M��d�sfN�g�$�dt&�D$j��`k�(QD����,�o�ߺ��������Ru��(�ͮ?��U������=��ϻh����K��푟=���p�<�me�T��j}Q�8eAC
[�)7���j�(u���
4Ȳ&XQ�߲�[�Ħ<���Ñ*�;f�R��J5HJg:+���1z%�����RN�"���C�r!���9�>1�Ӡ�7���H� �[[1�)񉜁���P��M��fQ��$4E�L62ʎ&c��"-����D����x���.�%+kd�����Ҕ���Ȝ � 廦�$@���k�V2�1Dč���ŏ�D(����I��km���VH㱥��6^I9��j.�@��ʱ�n�}��9G���2��瓀�g�����ݢy֮���ի��St�{.VD�G�`�@96�
$��ba`��UG̹������<c�ϴ_?a�9� y�����;��ƃri;�+%�+T��]a��_�\�4�B#^_g��*-~���ş����]���5
E�{^X~ֹ��ǨJ`XX�7�x��cjw�Z�JYNf��C���5	QK"t�.O�[�E�.]V�:As��w:,G@�ڷ��A4(`}iێ��[���am�Z�4ehf�S~����؂oM؈���k�r)��S��A�_�jS�Q"~���I�_��$N�Q-����=.�s��s��?����`��Ot�~�Gf��{%�Cv��^%2d�g[� j�sr<8Eu�}�zS�ݍ)�~�}Tz�£�8\� 4׿��XS8-�S�*Sd�?LX�@;Ēk)���KS.�Ekp�DH�5���t�ѡGe�O�M.�@�{��
.��[����������>��)7�{�n�3gB�Z�p-�U�׌zBE��P0k���С5o�S,Q ���$��N�-�)��<�ΐ�g�iJ�W�=;�uP���W����9h��],Ȅy5�O<��p��N8zq���lF?3���M���Q�X�|߾��rp?y�g��'��Cs��g���a�Sfӯ��6���c^W��>�������o�lL�鯾��[w�ƍ!/�<45��KVx)^�aku��[d�(������t�X����v�����4���fZ���j���!�Z��R��!�q�9uU6�I	�P $���ؼ�$�zn_����c�L��T���c �������?~Eء"���hk���7��0��u(��F��,�K�o�]'�xt��ˣ1���3:�����GͿ�ξ����zI�[�f�X��w�W9��9 km�$�q���E��ܯ�ж�%O��&�^�BH��¨�8n6�`0i��F��)�<BQ��Q˕'SM(�����j�55>o���<�a#D�����r�a��d��:^jN��]ĭq�������Ĕ� ����u�x&���c���^C�ZQM��K�y��@"�z9;w�<� ��J�7�����:��u�u����Sʃ���,�	���O���f�Z�X�B�<�Bɩx��v�*^�(�l��t^	01�����|��������׷ǘ`�[DD�l�tE�����ͼ��s5���p��ю��\wjwV7�^�_&�)�U��|DҞ\7H��Y�v��(�²H�G®��`m�I�I��	XM�HnB��~Y��K" n��!�p!�7km�`%�
7�<P�I<�6 �q�g��KFbA�D��	� ��W�u^�m�*7l�cz�,L � ��b_����9��"��i��Le�)Vy-i��fCY�Ƚ���E���(��J#��;�Ͼ�;���}X�=T2\2g�X~�1[+bn��7�m��֊�0�1g�5�_QJ�$���2I��X�������MyL�EӮ��J�
y�����l$���U�@%D��$eȺĳ�m~"��ęH�'�Pt��Ƹ������#����`	�G���D{~y��R���r��1�R"�v�����l5��-S�&�B@�:���bsB�J>Oy���YQ�~����laXR,�~�	_���.�㤥M��`eH�����s��9ҤP0�=���W'�t�&t����Aqe��D쳈gG���d-y�?S��A��F�Ӽ8���A�����3�e�L_-�NL<���Sj�ΐ'$�< 8��0C�e)7�>�p��s'�C���yC�f�q/m����P3�`�[=�a�Jޚ�yA {��"���#aË[CV�u��E��h��`g`f��'��VJ��I�SL�ō%�nX��+��"���߷6HZ� hY��X����J�(FN��m� ��Y��㿗���&�;9o��f*��/���9]��� �7~u�q�o��;�^z��M8� B��&Q)�]�U^�U������<g/�y�+@٢�J��%���RM���!u��^Й���RN��a�$��\h�
y)k��t��K��Fd|Z���>cN�tr��`j<ֱ��#[,���U��c5�%���h#B�|�3Ye�
X�:���D��1�$#B��!׷C�@!�Ʃ'�u�+�D�PU�L&��9�-bU�dZޘ�w�<� ^��膝����0���ʥJ�ZR|��L$Ce!I;���;X_8�-}����?�����qｂ7 'Y�X�8	���D�(���"X�Na�����N!b��~j��Ya�w��b�{���x���ͳe��=5˪��14� .�����ʜd�1ZQyr��X���`:O�?�;����[���1k.$���)I%z���g���ZD[ �1&8G�GN��Xۉ~�Vwwvs�{�u�G������]r�#:��	lu������n�5�kT	�R���;,^$ɭ�D�=IO�r�$ti(���m�H���� k0&�KZ$�ڑ�n��$/˒�'���vx���"@Wrc�sK�4|'���̫��y��&\v��a��N�!��Ƭ<T�ү�?PhY�Y,0& �\D0��?���������M�J;�I9s�,n59N������u B�{�z��[�H^���#�!�H䰰0��b���2o�ir��X�O��z� =5t�a�ͳ�גhB�M�+���$Λ<b��t���5�-o�� �ڤ�ȅ�1���Z�
�g<V@�5+rNQ��]�P�10iX��f���e�@�Ɉ�����B8�Y�fK+/1�/�56$�s�L(8���X{�^m�1�ڴJ�T�g�*Va3�y�^f�x�@ԭ������\�Z�)�jΆ}m�饯��5oz����;T���[���w��h�HJO�3ՔL��(�I>��秷��o��O�'���|.��ٺ��Um��� kL��*`�X�W�=��Y��&8 ��,5�zf���/\~��0���&���Ӕ:H��i�f}!���Y�F��GD$�'x���w�9	��h%:y�6_�j�1� �J$ͼo7[�c>� �{2$yRUA�2��'C��M9��Td"S�Lt���WI�y�yz��<�$��9z�a�^r�Y7^{Ί�Ɔ~�k�:`��S��{�p�;
"�X�v�uJ��R��R�Nd����$�1R����P���a�qs�?�)��J5��(aކ�?ޛYB���*���ߔ��P��o[����7�X"R�>nt"kEƤ�`T�I��&�Y��#�P�����s�������'7IYک�oa���Q���N ��������7����V��/�>D8���,O�s������A0�y��(�N#V�X1���[O�V�X{���9S�Yr����b��Gh�ZX��oy让	�~-4b�SnS�B^"��J�ލ�(�`�(<��~Q�re(�q�r��}��"3F1�i�d�Z�l��-��Uˀ���b�/m�0`E]JsI��ž������_uyX~x�<W��Ea*(Zi��.������a�\1��}9>w����R��i�Ӹ	�!�)-���x��z�kJ�ĀD�#�PS��/f3Q,�v���蕽�1G��_@��'���_��Z�X����_����J��O�~�Ì�_�O�|/F[���ZF�������Nd�����}p��o�o_���>���y��G�z��V]3��烟���o*�n������c���ť�lj1k������C[��p�6\zKN�V��k-���061XmL�5�K����SfU��JĆ?��	�/�0��M���'�;q���n~,n-�$2|����^���>�t�����m*ohQ7���6�nV@̄�x�)(����(�i�h Vm�*̦�X��O���m���������X���	�X�����7������Xk�5+�	�5+�=��� X�$`��C�
��RnÖ����X���܉i�q�JHR!�>�	S�<Bg8�y�ey�燵g��ζG�P=�f���0�����/_W<�K��n6����_�M��	[���Ź ��ZC=�GL����Ɯ�c��!�\-Agʣ� u����,R!a���QQ��������vݫ�-#��!SL��\�26��h06��b�j���X�¼�*p[���޶����5{���޳f?�߱���X?��?�g�`��BV]4Ь��կ�A@q���nZ��9�T��,���3%\�o��u�!�����l%�'o����\�q���Åg�(��6���YN&�<x(�S;�5�^�eCO��΢Jf��_��]��\Q5qE�,t��S-�%�+91M<ꬿk�v��m����C�u����4z�}~���$`��d�`e]o!:B�b?�J�5��ȱ6V<I�O������(ߏ�J�+�#<V�b��W����{X�U�ˉ�1(�uq�6����6U��zY��kׅE49����o5���&Q��RZ���rN&���+#s�xQ���-qݷOnR{�.g�c��]rSؘ�1�U_vS��4�R�Ӽ�tb(��G���9rj���D�d�4fg�A�;���N�?�i2{>���~��)�:�N�"â���	W 	\<�n�l|���Z������_:P>���������?؝ˮ��Y�$��'��K��2��N�.,�&W 6�VJ�3,�f�,L���j�֞�d<	n0�����x�(���8iy�ԇ;,���Q��pL-w���sv}K��P�5Z1>�.d#��W�E������7��ڴC�����$���'�H���֫����B��~
�;���t�S%���5RSyo��Q5��B9�q3�3|-�3��X!/
f�$���gM)l,b�,���x�V�Fn�A(�r� X!�!Y�)��	iƥ�d�L򬇻��ݢ~�2�MAU��#�����o���;�`,�#L�i	À/.�cԄ@[���J(�(ø�����
7��@�+}�"��Q3^=��� VF����
�tR};�����	���1����kה�h��T�zm=|㔍���:�lq�?�z��GpZ�kB�I��h�`߳�٫ V��+]|;���.�����{�o[�t��+.x�g�|牛��&�gOp�u��;������g䱪��ƛ���Z� 7���w:�-T�����NG�0��B"�AH�ۀ��i>�� !�����p���a���Z~�ԡ>����K�d����l�V�d�K~fp�6���d�6Y��	�"� ��,ڝ�쿹��pǏ��yZ�D�QH����wӹ��c��[ӦlD6uk�4�{��ʞy�@MC��x��Tn𥩝��H�v/+5�`,[���IOz2>����1c--�+��4<��:6�Jҁ�+!��ʱ���X��x���9ֱk�F�1��*�pm(�J:D^d���H�c �L�HZ��l���W�S��MkXɟ:�ټ1��݃�9�}��=+��3�ٹ�E�{��]��+l�5��@���Ɩ�([2��<���9Vk��5���5B���6A*'՟7�;�����'��s�����0cY�53ẽ?,�:
Ɂ�nM�R�7^���k>����N���q�|�H�0��ێ_z��_x��k<7�;[�c�\���ܰc`��L��QY����0����y3G��꒠!��Ax|4e���̈nW�UL	��Y�LYX�`��K�Fw6���ǈYOt!��<vZ��ӊv���\���&��\��a�&�� H�֨M�
ui��g%N�Y���D$��19���o�$ܰ�^�8��/+��Jm*u�թ^�q����|1J3'�E*�8�,r0��ҫQV��~9�xW�����S=�X(�4���&���m����~o2+䥔cų뱦P0eF�	��\�:��)\��`"?��MxD>�y^�ү9�gq�ᡏ��d)Q�i#xق���>uM8n�ju����w�`ɖ���8Rpz6�~��Ԑ��S|.l�=��_6lSw���z�	`�u�DٗvNP�m���τF��?Z�p���2/����0B��^J�Qx��f=�*�4���8��֜އ�_�@}.O����q�.6ä6�ݱ�)����˾B;J�CQ�8�y�����!�Q�*-˔h�;�TL��WЍ0�K��r���_%?H9#��Q_E[G�_�	;%A�l;�~|��Z��٦؄�ƑXlki-���m}��5�|�SW}��#z��ɐ�joI��u������5�}aq�Y�B4���ã�I��Z
�M�^��d��c���;�s�Q�����[�OI�I�*�-��K;��>��[ޫ��3m�]�H�Ɗݫ�[�������'�8]��e$��j�s����?������Z(���I��	[?��@)�ﵲ6����G���S��g���U�AM�ikƫK!�d�:�(pE���Us�n�.>��f��G|�q%oT��֒�J(˙�S�W�I�����C�E)ާ���U��h��v�`�
�旅^�F�������N�L~����X	Sns V0�Z�
&z��jcڧQ(؀Uѣai
��TPW(�e�y�q�g����S�Mw*�R��q,z����1t� B)��c�q�h<���>�k8����6<�M�j�G/ZSU33Z�l�P�����X�5���������y��[l�6  �IDAT�������ɴ�%;�)�����d��MҺ.��x?��Vw���aŰ����&����&��ŭ���踍cڊ����qm�>���E:m�w{��b���n��:1QK���{¾q~t
�m�i#;oנ�����?�[�~����Wo��>uΚ��Q��f���Eב]�^�I-��
�6��	�\K�h�)W�?��9;�9��-�S}�{�&�øѨ��?y�ݤ���\���?>tʏx��{�.,�t,$/�P�xzv���Qu��i�ån
��0�V�4���}(�^,�G}1mڶY���[���X�\k�hN�4���n̲�� 
Q����
�`����Y�Um)�\L��I��K���ևB��<�
�)�|M�5R�0���Ϲ���L��C@H��)���gi#��׮�/�Lz�5y�I���j�L%x��#ܒߣԆ<P������4��E�A �mI^�������gP���]u�<�# �AV�6R�;�E�F�&nb�V�4�m�q����ױJ~���J�F�CN�g�%�h�C��Ek���D��Ђ�'����fB=uѵ����K��r��3.X
>N�@UT(-b<G:�QU@�#��oC��jV�f�X	#3l�*F��>�}8��/�]ذEeD ��l�A����x�$1~X�
.�o���#�b�ᣗ,���|��5s^8��izgo�;0���ڜ�&r��G7-��m�ܰq��Y���Q���h*P�vn>13�܄�<��x��V#�)X���`N�cy��/jVU��S���LߗIAh��ۀc�[w�;��l�!�n�?i��+�[�S�K7���o5Qg��?�*��M����@
����?�Dʩf>1��WO>pc�4��k��Mm?��g߸k~/����h�V۸�b����l�#$#�Z�25;���|4iؾ��qӋ�I�i��2���I��]s����N�b�t�Mձfs�ѤӒx Ƚ$���9r�Q�_�fӅ�����x��BAV>VP�4����Z�m�J���mY5PdI��sD�}����W����cǮ�k�.�8MUGaQ��$�RU4,�~4�tc:u=��������Xu�~v�;"�FB\݅=�H������Җ���Z32_%���?����6�N�U�J�鳥9o���9?cn#0��&�Ph����)������{{�����ڏ]����2��ڬ��{=Xw�u�t��n�;��o��%��놏:;��햢��
�b�Ǽ�U�&�]ug� 6�E�b�b5�r�c��U���k=����HxՎ(g�<5�HlG����w�z4c�Q>cLJ��C���n�a��{?P���D�%�-�=,V�#k6�y��n��<���M�W����|�w�|��H�ڨ�L�$�y�#l�UV��I͡�~�L'�trx���-PL��T{��G�/��b��j������a�к�{��t�C7z�Q+Xq"�5Y3?�Է�3�8�D��@��[�~}ؽK,w���D�&E����8,	Xa���z4��]Ir���fŊ��|�B���������W��j��D�pӕh�]�`�XUn��)es������?/�;�d�<�Ϥ��he�V��	C��ȤG6l��E�H�s�O�7��PXϏCN�^r�� H9�Tמ�HN�`d��P���� FJGkk�4��ݜ��٧���������2=X��~^�;�� +��qc��K?������G>��>�|��wU:à�8G��.�����U5���Ѝ�Ny�h�Ф���g����Y�ڄ��Dڗ��6r��̘:]��62L��� �/�)��T�r2��[����jc��P�J7��N�Z�t�V��Xo�?}�7°`L�V 㵘JiH	�u�*��Y�"ʓ�Y{�����4t�I�o��p�I)f�~��뷆��S�' l����^��NM��Ⱦ�>��-�Kr���\zD�袋�3����lGWwx�'���'��Q_�(J��9y�9+�;3�%dwɣ�(
�-jE��w���T�t$;�Vl�޽��[o�V��:��1�G$�2�&�U�����3`��x�a�~�#a�fP�ڎ�0m	S(_�Y�-hI� ��p`��վ�T*HF��%5����)���͐��M\�ꭚ3�k�L5����/�;������*�۾eNK������O_v����{}��飼�w�V.L^_�_���)���?ز�om�aK���kP5eՈ���"K�^
mzWԛ�"�L.�$˞��G.���C�%bj>tZj�]�C59W}�ˆ|��!Q��Y"5�������V����[�{s3��k5�v+��t�	;��w�ج��������0ֲ��I�N--�c��n`ݧfy�KG�`���_�k��5�Y���G,
�<���/\�Y~�Z��zH��*V��b�c��^���5�h/�1�.+�7�ȣ��/�����!�sؼ����n������l�m<VB���X�^-�{��8�yy�������t^���۫s[��/���ɟx��ejF��k��l�4�X�tȀu8�i)�+.��z���J;�jYm�z���� ��+��+�<�)qX�j�c$�x������b���f�I!y��z7�iX �&脣Aܡf%*��n�p��Y7\��7��c���� ż�F��5�o(�rB��n~��%7�v��Ͼ���B����s�L.,������
g�)�r��.�Ac�v�gZ�k}߹g�_~N��7�dIg�hyZ�S�ҟ8q�7"N�JM��:\�҈59w�kr�Ui�7_�M�%��)_T�e?��JF�.��5p�Y��r�����0�L�(�q�:�c#�;���y���#R��0�~�>q��Êc��#�@Sز��p��_	�w���+W�E�[��A۸���4�kM���ޡPp��bZ���x�}�v�i��SO �O5�ߴ1��uכ����'>���
X��z�ܬP�[��tu+�|��cêU���,�W���o�=ܧ�섉������m�����X�
n)*�j���|�T(|��l��k�o_����%�:��;9�#L>�ܵ�ŇO-��^fd+[?_���2
T�yzO��׾�ݲ�Z�1��r�rD�
v�aX�ze��P�����Y.�Z˃����K׮[{�E'-m�Z��}|����k��w?�g��n��Ol���\�}E���o+����?O~RV$�/Z ���&�u3P�HžA���83|�K�{޾��YGeMw+�d��VF����C*�����LL�P3q�Լ�i�S&�7�s���~T�KɃ)�@Ɗ9�j}�O����S/����;�&��/�NՖJ9���%��Mk��/(x�j�+gG�v���R�PP�x��ma���a����|�F�}�W렶W�X�X��6¹�ٶ�lԩ��V �1+��@k�#��'̇g��`��O<��̬;���l����cXg�:�
&R��٭c��QLWo�n����χ�^���N�\�&�m����-:y�y�fX+]e�e��|�|��S�;�<�N��q��Vf��*Q*r8f ��������씧zWx�ɍ��k�<X���q��=I��
��N1��o�o>�S*CZyht�J�{~�����Xw׹MM𡦷C��i�����\�������~�#�s�H�ԃz���4���%(KG��I,B����[~ļp�ek����j!$��m�W�i��c�� *P���}2�^5�\̮}���?�r��΁r�9�،�԰\$'ked��B�b�J�s5�:� �u���C�rI5��K�N��0ʱ��y�S8�v�-ʥ6�Tlph8��"VOS��,]b���a�l�KK�OU#!7g�k+�6
ٶ��R�ӡ�n��4�҃j^M蕐-}4g)�<�g�q
:���x�XM$_![L����_"[��S-+bT��Ô�>d(��-�vX�ιs瘇
��гwy�o*�zX��>���Z�8c4t�jQ9ҷ7����p�/������>���l�J�#J�j �����uz��-�{�=����g��D���pe|�ێ�/u|	���fv��Q�����|���^��������>�/�M�<
yzm�Y��	w����}��+d��@� ��
� H�2�Yu(((����ө��Lͪ�;r^O�T�X�?gu���%W�wk�d�=X��=H��,z?+'�������7ޡ\LI�p�o�-��h�#zd��I�~����_d2�ϵ�:�
>xl۷���x�f�)�)�U�ک�	X�5`�qe��ԟ�Y�^�ab�:!�Vg����a1�E�+*��C9K�۴ȵ���kQ+�n��;U�M�6Q��yQݠZE2j��F�a��XƂ��:�r�X����nձԀ*򝝪5�����֚p�p}�=��Wظ]�<�F4�����f�����d�4��Ln4�y�I�s\8�;���w���8-9_��z�Q��@���ID0U����"H���|4l��rh��5��ч"��K�����[MJ�VϹ�.��6�
}���i-߲�g_����+�j�b���ˡt�t�jC�\nV����|s�'zs�k�XVnSK[�,sP&]V�"؏�l��I�J���,�I���:O��'��I�b�rNq�ʔ,_�>�զN���u�<�G����O�S�<��G\Ia#¿���~*��XӠj�����6 �P�UpW)1�Xԉ�kVk� 0K��4R�'k릟��8|@�/f�R����A�Pͫ�Ѳjc[
{B�4g��_�et ���>�j�Y��S�,'	IG��"F�V>��k��Ц�0�UJ�`���(�ô��ܣ�I�@x#���cͩ��P�w���8�v]H��<8��p_���^�4��jy8���ú�,M�4�3��߰~���9~��'�cOn�>#��<q��Qg�R=�bw�u]4���
��� i)V,�}yɬ�o_��w}�sNE�}�>ߡ)���xSkz4?~z����m�6l�y�@1�h�1;kjM�/+��h���TV�;���ʾ�՚�a���>/�<�hM�Ua�sC�\����������2�����x���sM�M[�!��.ƚ���Y��zu�FB��C�P���B��M^k{�_jF��-2
[,l밁��|0@ÛPПR�7&7S�ڱ�	��ڟ
��گD7�V�B`8J�* s�v��(3�3�Z����8	��Qc�<a��cXb1�/�:��}����_s���Ve��+6����,�l�y���Gi ���{����2�K��V�U�~XX�p^8��a���aN���;T����'�����%���/�^ںU�;���knM�x�qj�v�1�=*`���#My�RV1�yɢY�������Gm>؊u���x+_��X��H!~����q����l�-���dv�I��>y��� y;#�,ɭ�:WH�,�%a��R�9|��p�1��f��1�ؔ��I�3���v��[��
_�6��5�h���m����g½LyI�y�L�#�Փ��[y M����u�a�~K��"9�:�'��T�r�Y�M��%�Jh��Y*���h��ޞU��Z��STa㬑�%��P��:�%���3��N��/jC��|~C��W���sůk�L�D)��6Ā��R�'g_�V�����e�V�I��`�m��a���MpfgK��r�e��F�/#�0�m�i�@v��&�\���fTaoԫr�ۤm�
�g���K$���5���G���C���:!?�T(��{�:eՒ�w���o=w��}S���u�oz`��]n���������'�%����6{H�M��j	�@j�&*/i���؍��N�=9��SPr�3kA�� HR�G,��v�,���Ŋ�ЌD�<�&8�M����ԫ����06�~ �V��N�v:�z�����(��B�0�	�"��*TKad ��:�8�5��թ�~�����y��d|������K�hh�-+�L�	B}6�A��p��	beKo����,$� ��4�M\���2�M_!ǚ���l��ˋ���5�`+�ޢ�[^aki0�dB�[�X����%y�x�%��IG���/��4��O)���!�&�B�*�t,����*��B�ͺ�V�<4� �K��]�v���u�1o^�M����܁��Fp�����߸�Onڶﲎ�sg��|��Y�;�1�,�$:<*)[�`�R��	l	%&�&���.�#E3v���%@��5i36Z��Ǳz��TS��Ɔ�&��K�=."Z�ӯ�D��?�.�)t#L�%�r��F���kS��ɉ ���"@�" ����$͉�c3[Xi"�cڀ� K�b�i�����Il�h@h�q��A�P
p�&�)��8�P��&Ԟ00�sN�s�@���5K��s�̬��º�o����&���wIE,��G��R��*���׀�js�1��8əb(4�v��Q�&���j�l�2�*%B3�E���=�ݖ���w���O��CӠ:�����[X��߻q`�?�÷���S�^]옹RVy�71��R��I�(gm�`;�q���^.ک���w��U��o ��{��9��7[4 ;h?��Z���j���o�W�,zOw'@�~=T+�H!I��g�6	�P
�Ъ�C��J��ܪ�0B�DO ���R�j����8z�%+U��S�t��XSJśx��BM�f5���)9 +^d���0K]�3����#���Ds2�I �VI�i�&����O��̡z��п�c����h��'˅�^POkeo��&��z�#!�{��y�Þ�QiV�Ҍ*�����3�w�o��g����N�0}�܁��r��I����~rΝ���R��3G��;5��Z,�GW�E�,w:~����
L�@�`(ebW
Rv�Y;+�j̲e�;��j�v��|�!c-t��,J-�1�톑X�&n�%�g6Z��T�[㩲�i��z��E�E��)�f�Y�LD�Z՟?83��XM D`�_@�hײz��0�R	����:�E���weI��Cs�C���r�P����PmV_�yMŦQ�4�3&U��'�
�ց̣3t�q,��ƶ���D޴$Z�/J�мP��sTW�_���y#�Q2,Ke���l�?��m��"��>j�	~E�ԛ�)etͭ-BRy������Gh�nEp:���Q��g ݡɫzԉ���c�P��YȐ4�ۦ�E�s�y�D��$7<T�7{V~���Kf͸����t�;�yfI������[X� �_����o�Ƀg	��l��xT�fk��ˮKS^i��k�Z�w��RK����Œr��n2��(�T�:Al�Ԕ3BE�<��^Ғ^���~�?�YkkJ�v�V�+ce٫nHK\�����~��2�m!�Y�8��;h��{��[�;�>�"��)��G<��9M��m�	^���U�_=�����{f�bT��㱟!q��_q���g;.�g��d�΅�hpR�ap���q��XM�j�Hd��>#`,��N��� �qj�x���)Yy��f���h���3�a_��edb4�I��h&�G��֩����-\�]�G���2�d��q�m9��wK� �´r�����Fp��c�s(�9�N�7��.�ͥ)�*���Ӝ%Ќ^�&BsI/��nN^g.��I�3Խ�p�b+bc��ƎgV�^�Xt��M�D��%&���&��Y\�͝�{vm�u�e�_��+�va�5��}=W���޲�:~�HJ�Ltmi��]@k��^�y���6y�2�?p�s�{u����y&���D��j�{��zxM@���|t���]�w=�Fc�Ѹ�ƾ��ޗW
h{���*>��8���x��J�ѫ�����܁�k���ܮ�˘��w`�L߁�;��;0��#d�L߁�;0}���A��A@���     IEND�B`�PK   ��8Z�=�:��  � /   images/a3896090-6cd9-4aa0-adce-88a16a68907f.png��SLӯ�_� 	��	����;.�����!������������/��?LUW�\���S��"��A������ /���?���gl��@�� -����-=gΛ�)��Z�� D��!3A�F�kHv������� �s���1Cר���ސ��)�
��0�L�M �~��Sxx�-�[���0��1�:�4�Lr�<��'�K"@ $Iq ��\1A|�?jf��uѹ�#�� B���
��%����&��ڡ�x>@"�/��J#�@�_��>�ՒV��?3�����-�
"��>��D�v��/�_����B�����/�_���аW=�����,y�����K�ǫ�3���뮀�n�?ۜ>g�T�s���?u�jQF�dHO�aOüthO7b�b�HmE�����τS^-骚��u�i3c�/M��K��Y�(F-/`�Fݏ�	�7{_߽�a@��Xک������)��/�i�z	3���*�̉����(��u�{rq��YԷ��O3�D��Nɞ<�5��Y4�6��/�P>;�����N�컱oW��T0�v��g�����63��V����	��z��Z�JL��z��X����i�5Hp����y�G����z���`�w�����t��~Ԍ�zT��Y/��\?����J�8���3Kfd|<��Ԉq���:�r�=@�]�^	�Q�R��x�U���LB�g>�VQ6���?�:͚����0�t;aQ	���<�6��D��F�ſ�|'H�0��^s�|j�V#A��.���A�OoK���
��	������`��JL�-�)��1Q� j����4Hׅ�أ5͉�1H�m���-683_@P'ژ�s��F7Q�'j���a\6�ަ�9<�����O߭�8�%��z�{�Id?�ф������=]��EXg�K>�+g����H輦U��>H��;F.����c�U��{Y�t4Ä��A`�P���הզ��%{� �[F���9?�a�9ѻQ��*��s�YU$���̟.�x��9���ԓ���布��*����`�^v����tϷ���ߒ�p�ru��G@�'�V��dW I��O�t<:��Īȫ�Z����GӶ��횄�{�{�\M'ų�+Bh�TBTl Џ��k�%@&��e��v�m�g�������$[h�A7��>��>��~1=U|/���w���j��z ©�u�KX���W*
���2*4W�s�;�.�]o���څŬ����ۆ�w�)2z��>��/O��[��u�����5> �=|F���n��?���w>��R��	�֡�fWΥc+��t})1E8]�����*�Y}�f�(W�#2�'����=�w���Z���(��n K���YU�X!�&:���w���/5�e��	�r[Sv��h��΄ef�K�C�xS(?E�I8�x�D�SMҝ9�(��$m�h2�b� DH�L�A�fn�8�쩕�r_�.8&_i� (�?��ca�Ι�B�G���*�~߸c���a��D]$�j���a�N�0U�#��k!���%�|�Nw2I#'U�E�L����X������>�[����<�_�ހ�+l�޲�L�PP��ﲊ�Ez����,��]�ϒ��/�fP˟��C�vqy4�q�E?rT�V�:e���Eܗ5�C_.��ôh��pO^�hn<U+�)+��$�n�ט��0`*g���в~h&�ؤm��k����6Z��	ŃYh�QJ\,��؊�����#��������Oƙ��7mբ���޾��͝�m��.���Put�/����b�4{q�������@C�+1&�����T�b��^�%,��� ���2�돽�A�f$�J81���vs��_;/�B��)�e��qQ�<�מ]�l���F��M�23�g����#ޝVsz�I@�F�O�3X��	���o���'W��?��h�]� ����/%�6�W2	�����W��g4Ŧ�bɱT���G�(��Z4�jф���:�����Ϩ��2���X�8$.����5��GzhY	C���_�'����̻�ic�!��-���8ct�8[���Ʉ�j��%-�����{��hj�sav������+*ٶ <g�`6Tj\�O�Ɨ�^�_�����糪/��b>��J݌4Ht��-b���f,Eo�1�_<��O'1�cp�X�)Icp\��zF�� j���Z=q�9P��ؒ�V=�3&
à�d=�'i�]�^]5�+�It���^�)~8j���(@ek�� ��Q�и3̄�&[oV,d3-���Jy��%��b��J�˘�)|��DA��_D���3�!jNolvL�d!%I잫�պ���)z)�������/��W�|\���2}aH<�K,IY�Z:sX(=>���ZJ�HΣ`$��QJ_���BNl2��/��R�΄İ��򶏏[�fw�dR�g���s��&��?��Np���aS�����Fގ<1;��{!�f�c�8���P8��h��΋Y�΋,�I;����#�F�e�����݋%t���V��'9'@ǌо�M�����8���2pg�	�f�����˼�r�V?W(����r2�����5�(c�0�G>����BfN�m��J�0�Y�)ϫ͘�J�\�,AA�܄ʐ��1*𖌖�jܚK-p�����[�H�-�Іh��W
����?X:�����Q(��#�=�?��ܟ�����^�lr�r	N�6ER��	&���
����D?�m�K|�BfDw= ����6W���kk�l̶�;W��{<5�>q8h��A�lg=��Ƞ���!-Ni^�`{^�a.�^���써�eR�?x�&	���遘�}��$%Z��|��d8���/4�2b�����J!�k�iZt���ŕ�f����e��6��	 9����h@W��W-Trܣ��;���&}!k��� ��ݻ{�$�}TX#6v<�%������-&�Ĺh��Oo� xN��L���K�'ں�u�^w8Y��*;Ћ�����n�&���U���ݦ�z�����ݓ'?߫_��&�;��>-�x}�3��T��d�(5$�J2���ǁ�Ūŕ0`֎,�r,�����1�*
[���I����t����c{��3>�����b��|��M���&C�ʬ]k�i34��sPٟ��&ڪ��_j-�ץ�1�*>y�_�RɌ�ILD�d�#��f����4�0j�4勧BJ��!gF	��`���ڿ�4�-ؖ�% �ذ=n��W^A�#�}�6��X��\��4#�?i(���L�
�~t�.v��Al�[� X£_�����=��"� ��ݓ��4'U�L�Y�s�-�(ne���}k!��>�HU�gT΢u��p�{�g���#���Q�/��"�!����˪�y�лh�:�������:U���x0o��D��YO�.�y��";��El�ݤ�6��.�ߦOV��~ڞ��$��_�����4-?��W݇�e �a�kK�k�!�8用���==���t�ʶ���đǇ;Is�&z��D=��Oeq� �_�wrG����պ�U���Ⱦ���> �!�2�m�j<�T�麯����8ꪈ8��x\���vß+\;���6��^�2p�;v���R~��tGjs�1?"O��?i.+�$��/��
q����|ӳn{���ܘĿ�l	;��Y�d�B�6 �������$��<s���(Y�!�{�G$ (д����O��Q��d�|���)B���X�8��,����;�V�����یD<]~��DFGB�/�,J�O.�j)�gWWQu��^)
�4�sO����`�\�'�\�cZ?*���9֐������+�f����nGJ�㓲�4��Ƞ�,��֚[��8�>(sΎC�� ��|N��s�X��8ט4�ý�A��G����,(�x�y?\�	�-��~,Es��S�	7�S�{'j�#�8
�'�$D��D4]�	!�'(Ԧp��a@W{c����C�{H3�@{�׸���	��Xp9��k�Y�Й/��E��� N�A��ʪ}�&foZ�=�ȉCЕ�*� ���elsC��C%bXp
�\�Y����xr�"���6�93aq�F�7T����5��ci��i���M��!�\���Ge��Wf�w��rH��#Y�?*$���%��gV�>�f*@{Y�9���ra욅�kg�v.e0��(���cC+�χ��"M�9ܷDZU|�o�[��uw����M:`��@rM����;f�ٯ&%���i(͆�v�/�� ��n���bL?��������5�~�R�"d� s��ItX����D�6,�Pf�3�9	ʽ���i�\<��췖�=�lr]�(ڷ/�<�g[�/������4�r1�U6�n�%���͓��(4,x۴"T�i߾�l����b�h�l�hN�!��4�MKƶ��d�SNWO�x.���H�z�-p����+�\JұҺь�=}��!=Zcr�x�7����ے����"P�b�^<<�ӡ�mKw�f���Iѣ�Y��s^3�]���������S������������%��q�p�bg5l�C�n��~(�x�5膙����<h���ߎ�R��b�GQǡ�'rJ&A�r{rE�&|7��(0~"�G��V*B�S+�]]'ܸ���ZK-�	l&���wnhE���q:hҢ��ȶ�оXL��$��Y���D��ϡOQ�
 ��]�V�A�&Ɩ=�y�����w�ƒ���o�upy��N���[2��i
I���7kQ��Uf�tl�Ȓ�GS sP��:���ᆧ,G >�Bz����� ur�.˭o�m
���������U�V��jӽ0� ����G��<��|MV�񰣈��m+��=��A�G���&T��ʦ���R#�4??�����ǁ��M�wn���N=�Y$���6$X�js�C�c�ޠ�\��~�|�	58��+G������;
3��D�Q�36����h���vQ$�H�=cA�7l}��:�#���^���oШ�h�+��IǴ�,,���U^޸��<���H�au����P�]�m3!8S��V�#"����'��.�u�
ƫ'���TZn���q秪���D�dܻz6�P��t�BK�rHGzp$�tXjH/��I�W �	!�S�E����`�OG02e^M잯9C)h�%�K�1��í�����E���+����OW�MTV��<���h:h<�^�������}�h@����]�(��3�I
��?��+%ǵh+�O���>:=����|�
z?�1S#�W��>|��DR��,��	�9ol��	�x�I��ѝrG�TK�t�a���4���s,��p-ӣ�6�O�P.b���a{Ӯ�?�����⽟m��2��.(��~f���^&-�����H+�g�	_�N%��=�����>�l�u�|���s8s�U�._���@�A��踙ҏ
�֋n�nS�]q���1���I�D<A x�ß$=ς�����(Q��w�]6]CI��FHw�mu��F�Qf���]���Xƃh;��ˌ��B�4�>�(bRT&[�n����~��l߱?Nl%C��"-��%B��W��>�4����hC{?
���vNh���f|�1Ν��k9*:�GЉ�w>O�y���7Ѹ�1k��ﷅ��6�3�GKT����t�[;�7�9B�Ý�/Q���X�~���[6���m�3�FOEv'0j��=6?���b���]��C� �&5HYo��i�86��SB��|�Bl�^��Z_�)#��4���W�����:���w0?gە�<7+9ɒ:WC�)���J~dDW�!!��I�7���T�d����ic!�R����R@�.ɬ�2N��S�э�#���k<�H�ʝ�~9�f�
��Vi`5t)Wv	��&�-0�!m��:�)Z �z���-:��)*��LI�,-����[�5�Z�o��懑���N�8a�Y�啼6N�^�.?�AZo<~�	�T�>��S�����y+�'�z H��$�����2�A(�J!Zz�:)U�~�!����}�Њ�a��
�z�@IIyڊ�q�k���o��0�j|j��:w�旺+�V�mLM2�BJPu���q�a�݈kv�2}L[:�뾻�>%!��$D�#y,�̶N�@W�?���}���<�.9����m�-��C^�)2�u���4G~�Nxv�+��83{ ��F��D� Q݄��(�2�'X�I�+���6�w��D"P���{e�K� ��Pd����w�����t~��G�x@0M�x*��o��ܪ�� �x�T�����N��=�]�L:���wE�k�o���Î�&0�bl����{ V�z;4����=�
����F�q�������pon=�ۮ�l_f�+8R;��J/}��/��<����*�_7&ײc>��Y1%1
5�����j[�a����g�PKMߤ�`EOޛ�² fs��ZC)���D	2�b��T�Z������+���Ϝ�ǭ��FP�of6{7�dgpۏ��C�69<�1'k�r�#�A�'�1'O�*}k���+���ÙƾȦF�&V!�c�;k�o42������pH���������Ӳ��+���2��^cE֦:sT�}B���H��YW�3�I:##�P��0����yf�Hh�ŵ�uĆ��&�gz�W�H�Y���e�[��"�"��$�}OCi�<4:]�փO]Ĩ�	-��Ct�Ro+鞨F��޾K�R�gp�gPh��m��
�rK��� PU���GS����{'��6nw�C��w��@|��cE_狐�����BŪ�r:��R!�S��g���7<�q�F�:�z�y�yrL��k���4^}����v����V�$��B=�-}�FHpj%d�Z��o��k��̱P�fl#%ڕ���,�mZ��6��V6���W�H��<�!��_�>��5�;܅�T�AL�x�����.M$6�ӼK��b�]-WZڹN
/�&���p�*�h��Q��/6�sj�s�AlUK�|�C�E�+�)�Z4��Z�m@�[��N���F�๟3�O���ύ����'��
�3�1���y�gU�έe^�9����0E��,�㇉������U��Q3,�B�ږ�͔�!� ����" _���̒��hf���
��)V��K��Ѩ��/Y��!!������JL��pM����o�����[���v�ڿJ��'m��?	1�܀�� Q	��V�v���������S�&�&�dh�8�(����{ЮRpZU�7S�ɗn��^G�;��%%<��4�����;�GQ�C���:���7����"����-�^�#i5=�=�D�&�=&�0#�-�ԝAy�3��G�v1�`ƠﱑS?�B��=�ʗ�F��|/>E��r����c�Q'�k�+�'����xY�UC1z΋��z�e�\��6��%�i \����L���l��J���;*�n��1�/>vw�DA��>��3��}����x�����M�����ꟖŘ��FŇ4�~T�w���L���[8]��R�ͩǋp
V��d����b��Z�T6F���bnE�Θ��vi{1"��4,�������77czަ���:�(��w����%!G���vϕ��G4�\I6�Km( �l|��|Q@��*�[�B=�<�H��C?�_���s� �ɪ+����7����W��HW\�|��o&W7��Ksn7��<������I�h������s �h�儜a�G�
{,\�i��I}�0V��9{-[>��49�Td��*r�������r�S��fiW��h�IOܠk^�Ej�TV��E|B���v�z���	M��aQcꇞ](E�	Z�E)��Ê$�둞"�b��~u��7�9�=��e뚻=^�j`Tm>�n8)!wl���EyJј_�F��M��?ƍ� ��ZkM����I;���O�^�jN����b�?�����������Ȳ��e���t�nC��o����}��}b����S)��%%��V�l���
�c��+�m�������Ԣ��x�F3|��D�,�6.z��>ٟ���+0�[^�D^f��9�f���:|����Z.a��}�Bc*HN�X� ;QH˃�gsˀH��hĶ��$h'a��U#��S6��)���������{������>�ؤs�u�%��	�/By�_<���w]�� ��-�2�Rlf��ws<�]�@d>1����w냌��q>����j}H�S��2�Ѩ�d(�1�lBǽ�8�������Y��%W��h��4Y��E����~�����j�s�R!=�F.������Ľ�*�U����)+�J���K�rF ֺ�IOZC�Ĕ��М�!Wȃ���i�j�K�@y�� %�N)/�b-��`1��ϔ>D�Gv�Fy�U&S��$��=��Oǫ8@��5�(|�s7��/晗�xU���H�g�i�6��4�tS0_U������Tg!h��m�Nn�a]d�/�Ƽ��#�~d(�6��l�z�;�N��q�ܪ8�4B��+$���>�����ޛH'��~<��g�:[��z0:��\e��u,�9O�0nCUV8��s�<��~4N���/&��r߰ �+҉�}P�u��L�yu�ݹ�;�W򬚺&~�N��<��.�"C���J��|Vjw�W:�~<�H�i�#-�Xn�����d�|Ģ �V,�}<"6�o&V��r�(��[{����v\�f�_g�پ�v�M�$��/�n>�e	�JJ-�C'��n��KάW�s�@3����\��@޵R)��r/��f�5��HL��%$t�*l(F@��|0������ވ�"��g7�Oo6�Ҋ���M����o8���&%F��Z�Z)��,�N׎�����V��"*B�� ui�lO�=�D���l��s�/�
�#������8��h��V&z>��9>^�Τ�l&{X���adg(�a;�:m��.l��S�K���(+��aU�#曚�u��*���>u1,	�A��H:��BX_���[���J�xi5���TSI�Ս��3�ˋ�,���t�vV�F�	Ni��X����G�?a��i*`=�� v50�,k���g%TWr{1����:��خ�>��M �h[��?��1R��!��	�VVwa�Y7u��Ň2���g�I��8�_G��#<���G��I�[��<�>��5��O�?�\A��q���Tsm�6�t��(�˥A��ډv����ӗ=�
'P2���_��8֨�6]�vRˆ[Ex.���~�ݡAn�+��84�SN���r��ޏׁ\��S�۷@"W��X�sO������<� ���_���� �����}�K@z�0��2��D
��sɼ�������dA�^�g���퍕.�ܯ~�
����TB�3@����kc�^�g'.��^5翽$����z5|����1���a���F�:i�؈¸�P�� 1��y������ia�.@5���f���H$�| n�E�6<�%}��8̩E<�E�]F�V8 �vX��� ��,aK[�I�8̴�d�h��b�$�%Hʄ�#���GT:�A���F�٥��;?-��*�C�8yw�ЏEh��n���[�_9����]$ (o��m��ן���J��e�S�x/��esW?r��8�Kw����Z��uQ�z,�=�z��a2Y*���5L�P�/����%I����o�՗bU�o�C���B�a4�%�u%gR�wxF�uqK�}/��iWϮt�E�rTӆ����8���
y���1
"u����D3M6�@$e-�8i�.��>�f��bh�x����r� �9a�l�����q�X �v�w;pud�Y�2�ڞ�L�p?stn��7!lߥlm_GO����Ӯ���e�:���FP��(�iZ���Q���J������&���о��d��2��}4����Dʴ�����nyE�ny3��ͻr]6SUV�q���nײ��@���\B�q�Bn@쨒5F©G)���rU3E�}��I$��5A��Y�ۻ����	~��&kFǔ
M�	�u�J9�ꃡ�/�E�gE3׉��S�Ύ��r�����8 ��_��r=*�G�fqr�Y���A��J	�.예#)����o�Cή-ǯiY���
�x㟴=���`�v�1P��_\㜍��pc�@����u���Bݩ_h�4��C-�-f�٣���E�����/Ȕ�ם��{��s�)ݻˣۭ+��e��N�H���?g��O���:k�d��)
�H!�}v���_��"/�m��J�U���Ju��~�q[��]����D-e�1�G�X�́�a�P�­*ߺ5�p��{�e6L�������͍�WjX��i�E���U��������d��5z�ӫ�e���vũ�S+5�Ϲ&��EエW/���󈔘�f��1{'��ɓ�V��t��^,~���-���Y�g���t�R������"R��9ꆅ�u뀇X�޴m���R����S�bHB���c7:���_��{�q�:v��/���mc�����	6�ښ�ub�z�#r{.�{�M�`����_�?]�B�pN����n-���bGS�èv�b����BC��h9��-&ҍ�0j.�:�̨v#̼G:�:/��2������֍�#�(��35(1����x8{��/�F�e�� ��3��_�f"#a+]o�絸q��pm\��0�=e��[��.R̙)��u���%(�1Y,
�
Ο{�`G?*�1��i��S�q�����!D��7���P�;�X#5����ly46?m�"yǪC�r���ȸ�{|-`��b)A��A��¹$8�J�;���6b#�3��ݳmB�L`�5���cvNe�J���)�,�',MdP�˓j^#ai�}�Ŕ�
+ߚ�
��{u�e��T��-c�p�IPUc�
?�#�y��i:��DX�H�4�kz]r����Ylv�S����R����'WR���Z�Ĭ8��$�Z.5�V7Y���+	ިپp�=V�8?�ߦ����,7�-CU�.��@L��`}��Q��@���ղ�9}���o1�9�a�D��i�Ǎ���}i^d	���jZ��q�ÆR�m	�����ih�8�5�����2��Ғ59_�$�~'%l�D��6G��N*B�DZo?\U��j�y��P�yFl(c4Ŷ���A�|K��5A���Tf-���h4�YFl73SQEH��b��.����8���n���::�����#����8�v{1��O*eտ�-�,��4{����\�2=f(�n�-=��[��}�.�z]�coC*�²��gf��U<:0�Zt>�J�HSx������/�CUz>3�٤�K��������U��&(����ܳ�ran_e/Y��л�ee���i.����@
���ԼVg<[���_Cv�F��WC2��FsƏ ��֚di��fL
B����[]4���Řv�����v��3�p����=R��}��0�-�@���r�m%t-D�q�|};I�����Y��5׽�D��bS~��������0���\ߏd����Jiv[�$��O��.�_%u^�\Xȵ���v���o�k%���f�kj���ܞ��P��K[�"��7��k=gJܪs0�?�����}�RI�J$��m9Ƣ�c:y��>��6Qy8���0_1���k"6����-=,���'�����̵���D�����'�lqEzU��L�ȋ�hT��ut] 8V�P��0��c��!�I����pkf�K$N��6��VG�az*��Zg2�\Bey�nW�չ��C�GP���S�/f�}�.�����]��	V� h�T�R�je�2R�qϚ��zs}���V!3��_��!�(d:X��Z$�Y�!qC��$��a�+]�M��q�l'q:;�s�zm��0�Gf#WA�k�D\���w(TS����bY�c���=q����/wϺ����/�t��o?/Q�� �~��:a"��C����,0��t�`"���N�����xH��x'�},�4a����=�c�;p^�)�Z�jȁ���s�m��{��yi��������$�;�Z����};�$Zí��F/`��w/��	�]���;��"��;��0n|ؿ�
2=W6�;�6^	���v�@+�|�k����B~W?�ۚ��pW̑���~�r���]�}�v'���5��(����Y~A����,�'��S�~�ۉe>{�,?�As��)3dd�y�PQӣ��̯'�d5�sC>Yk��Gm�_��W�Q���l>�Ћ5y������Xq)�
5cR��z ̕��-qӑ)����Χc!���Z�q�jx�d4�Z�� �s��<r�����M#����8����0���+S��o�p��x��f�Ӿ*?����;�!�)Rw5�<����I��F����8�3�I更�ԍ�c�>���RD4{���Y<*Q���؆�ϣ��i�=�]�1��<e��wZ����N�ԫ͘M���r;���{�L���dG�����j�=`�T�����(��J�w���V��	�ج��b��Zݔ���RJk�so�|�	�R��l�Q�Ϣ���2��m>�c��,�Yi���Σ���4M��-Ǖ�2Ĺ�h�q;"��
�/��9k��^��7�R����� mR� 0�&�^�8��Nz,]��7 g�	*S��)s�P1��Y~�	��!��[�s�۽�30�$�wű)B[�7�Dc� �g�Q��C�:#g�GY���܄N8;�u�)�t�ہ:�E׵m�|�:5�'IN���@D@ �@�¹:��:�����n���o���zn T���:�s����c4�3����!3O0�%x�Y�Y�n_��>:>�l��������hZ�Q�y-�ah�
��t\v`���6ĵ� h�4%7�b�q�����\9�i_�X�I��kΩ�m��L�[����IX��0Bd���@����\n��<��J���[5{:��_�S�'�BH�@(���e�sSm�wē��%��@��q+���������a@dV����	�P* ���,v���0QOia�O".W+�j��,�R��+m8 N���8��G��xj&R��Z�܎B��S!,��"t����۝5�+/���+-�a��^���
'w	�[6�v��7��j,��L�r���h�2��S���ͽ�����W���ͦ��e���Y��)j>D ��&���c�/ �fm�2�%K��7�O������N��3�VF�>S����r�r���D����s튷3�p���1(�]6��6tQ{��H���7��w�"U"�U	)l}�T�ς��o�Ux Ch�eJ⠲{}q�X��)�Қ��ô>�֡o�u>�BX;{�ʏ�b�Ŷ�lGX3%�����!���DDs���!_t��Ɩ)�$Q��#�V��������b?��#��Lʥ�I�H�Y =���( �(�o����z���~�D�5�;��gB#��zDJa��(g�mϾ�	_�2�rC	z�㠕���/8�'��@M��\ĝ���*eu]�\ �M4씭$�լBz�M�[���0O8�;U�>���R���x�)�w<c��}@b��ot��y�÷4<fĞ�����g'�ˇ�'�b������4���D"�r*��	�W���1UU��},��AF��i%"oZ��)u�;+�����/'���h�	����L���~��Z�����Fn�� m8�~Ӊn�w�)"��\�-p)s���3W��}��/c,�#�@"�v�X�b �O� ��Y�X6Dɬ��1�4�!�C��:L�R8ct�ęrH:~L��/�!��A��+{fV���C�/�v
�0�v�P�G ��4a�2b2��]��cQ��dϘ�fqN�pQ�; �G�mJ�K�W8�z��l##w��O���h�m�޹L���v$]�
[i3˵[q�9�h) E:���q;���аj�`u0�ϑ�Q0c \�������B'�B��X��D�}��~�dK���1�3TO9���ίB]5��7y���j[�A�~mY���S�� �����`�&�}�rOL�ӄ�U��#o�~E����U�f<5["��wɼ��l�N��0x����r6�#�yϖTK�׈�wy�'k[� H����@�Y�Xط����<�6OG��,��wUK;`���,�H��O2�OC(�]�{����/��mSc�<�lǻi��g�ő��w�&?�ɔ6�G���z�/��9��@SqޥM,��~-4��T�tGPj>��/���!>R[d4t�'�0ΰV��-�<4��;�4���z\D�����0�ż��'a�]z�t>�-I���m�E$��\	�����#O�2��C��,�/m]ix:�?3��B�#ތ����|n
�bf��BWyw�I6?�kS�1�F���e�D��N��W��t"�ҝvz��H�D������ż&����$akCz�*:�UԵ�y����D|&]�ƾ�%�X0gi7g�cə����w2sk+a�_1�gϻ
���T[�����)��^iCcb�{<]�1~%���pݎ��`x����٢16��=�j�w(�j�����+O��S'�
��v��,ũ�h�36��O�����2߉�:����	{��Ya��	���WQ�u�$W��C�@Ўl?M(�_#@��QC�
������e%s��L}x�J�q&,�wC��3�"�$�A�=�c�w�{;�]<Fz�O���-T�G�L�o蓨y^������R�=@Q��d��"�	���n�������b��A����ͭ�^��?*����!ԕ��xzH�"�� O�e��E�*0\"H�Fr�ׅ�Xx𧤊-&:o֢��w)�u�� ؋��dYP[b����[��Fg�"w�o�卟Z���r��~���%g��6�t�tɝ6�����UE�|oPM�\쿠_�~F�NwFB�V�^����{�����;R�jaf)^��o��i�7�7���ZqΟ�(��~#a���('B]�����*�a�����C0ӽ�L
�{����F���_*H-޼i�V�_����	Y52�S��:�w_HMLg+a� |M�oal�<Ze�6�"ۈ���	b�"j|�(%g/�ź��qL��|�
4J�O�gMW��㑫��(w�pZV'Į�(�On�j��+S=�4�P8�oC:��v9�,�}rf����g�.f�"Q����Yφ�Z�`��⻔T
��.7ň?�ȍZv}�k�����[�����ut4�A��|��ڂɾg'y�4����O�$��j���}�B�������6溧�c >�ؙmǗ���{�3����
� �Hҍ�'a�=�MQ���r�O�������hw�!����������W��Y'��1����5��-���"/�1�H�T�AW_f����\~�b�;{{G/sJA��Ѳ�M��1m�o�;�r���"��a�ZiM	��P���V��_{��iRب�1ծ$]�{�HZ	?_��T�a��rj�g���>��_���;��ƓO�in�I����]h��S��>�,b 6�Q͌�����Rׄ�����wx љ2����/�5����x��)+2��1�Q�C_P�݅�J�#����z�2�����Bi�:щ`��b�n�b�)��pJ��8�Ok"F�=RT�G��+*	��,JK��ܤ�%��W�Q�4����߿�#2-�"�]�ǎ{Ʊ\��F��^黲U	RpU�J�I�6��E34<�8d��t���p��FN����CWS�v�}�LdDc����j�[1m��u�qɘ_7*�W�U� �t-f'[�a��!��t(]��z;�Hn7�β%���B�w��P�=��H��2���Xr��ޥ�'g@��a�fd�Ǐ��{����@a���+�N\�2��6�䆍aֶۘcp�͏n5ŏ>W�E�)�c�q�k����`�j6��=p���W}�}JF7��s�����w���h��dzJ}�Τ���?�&�	��8�+��VҒ����Ť�j���d=�]\:�!�SC�(��[�du'Bw������EN<�Vn�:��
�OZ�j?�*�*ח���koG�l�\I8���E�q8�f����q��>�������e�|�m�k�}^p�M�Ext=޹-� � O��B`�����6��*�y��j&�"i�T������u5�X��������'��:
�+��?T�eS���ܭ�)�����xqww�k�wk��Z�xpwww������~;{>�sfO;�F�P�^�J�ז3���i�Y#�L;@���Mj���<3��ŉe���(�wB��C�.7)�ٔvh��~��~ґN*���x���ǻ�&���F=�"=�J�ԩOW��c����ET��ǅ4�-�yJ�N�#zM��5��Q���U\�G�g��5�1f��5�J��H<^�&j[�-��`Nx�}�/��R]�g/iNg�/��QP�L+`����
h�|\,��V�R�Z���7��-��:��!�oL�qC���
A�Տ�P���$�耰'}Y�)�a�2�^�GLy��Ü�OC����ʞbI��_����{Yɤu?����왙�������j�q��S����\.8��S��L���eY cr�E�ߣ��޶c���A��� .p�c�4�b�o5��Ҍj��ǹ�=/D3:8�-����>7o��i�����>Ӈ>��qU�@u���b�*�W1(�'��xyX{���;V^�K'E���PX'��Oʹv��\�V�F��˪��
Iy9T>��g]e�◄Z,�3ޜ���d�y=��F���D�	
۽?){#/3諎�_�K�"��%If�ܦ*.���7i��}�S�S���b��>�z{�=W9I��k��[�e�m��:�wT_�
�+��-z�h��\_���;�|.���z��~�$W
L���ܷ��g�s�lEt�gD$E�S�S�u��j���g�0G�@�M\ļ��P�;8I���{�'4�^�D���(Bo;�x&Ǿ��T�C���>��cq��_Ll*��鐞Tw�2.�X���0��KK�ν�J�'����p��V)sW�<x����?*9� 8�z<���xz5x�%��&r��4�YM�4|����;1�����7kY>�����f9�nu�vP�d���یI��Cg �Y��/]�p�#t�H���_�Ƚ;CF���S���u���ċ!���a2u�=f@"M��ElQ�Ւ���qWNq�FyȠ�x�O,�Ґ�'��p��v,4yu�X��[�kOK/���j���>��U�u��� ��vȩ������%	���s�����/~i�m��$A=G@�+�M:8҇;��;��m��1ư.a�<��Zx�)EkU�({�ﴀ>�<m�B��qÖ���P�v/R�33�K%�q�*�M*1|�����&x�3�yA�5J��'�e*ӛJ��<�Q���.&�|u��,�������-�ū.1��| *4�I�bC�%4��߄D��>�ߎ�z�^s�=_rJ��x�x�0u ����r��ㅀ�q�5��ĝ�����i�}p��=42�XF=����������
=u\���W�h�-s�:r�m������$���[�R��[�E�2�����O���
���q�*Id�Ձ;MN� ӫ�m�2�n��ǔo���A|"�NF���Z�⾽8@��cT�C��}��PE�Y��5���^���V�r@�(�%��^���ι��	���j;�:R�7��A�$9���c��ө��D��I�e$�i��uڻ�/!�oZ�X��\�����U1���jS=�F^0w廋�r�
cE̽��z��Ia��R��J�S���/����a��gq������B$��.~{TXu�M�`��Ê�>��;�\�L�tܔ3�7��"�g��`���6�v�k�Ð�5s3|[%�%K���_-�7-��u�e�{�9V��ٻ��LY�J�S��N-���m�C�1���Uw7�@�C���O�e?j����d��6�9Is�&1--��P~%����C�G.���L'LsGO+����5ƻ3S�j-�����=#����ﻲ����n������q�u��n�'�{\��$|}p��ߵ-��Opo�a���Zk���@�����	��I�d�ĞN���8�9�D�n�	9(:�����@Ӈ���%'l��ȧ��&�;�c���@��1���H��H�7#j�{�H3o%͑`���G�)���%�ѡ���T�;Ow���[ƺxI��o��`�J3O��
2r�����#��G��,u�����LgU�����.�X�{~4�Kw�Ґ:��C�%��V�3�j�5q��&��c+�Ƿy�q��$m�!Z\%���1����+u||����`���=0!��L{��&�l �k��𽰼ߎ�����K]�DW����3���e�����S5�l&r������¾����m׻�]�b���~���{\�o���W���(-}k���3��_�ܰ@��� Y�A0���aB�C�ނ쏱 ^{��&������������?��-���bq�������p':���|w�Fq� �8d,_�*����(;�\�b�hN��s;E�o�
�HFD@*}�=��	=�I:ُ��Mc�F��g#�$��*OCp��C��@e]�u���D�T sN���=�?���z�����O�KC���1��6�w2�a������]�L�O���D4���g+4R�h!�/�]�+�{��ryRA��GA���M��$^~#�0Kߔ��HX�N�j�:�P]Yo��9�K�����!|>O�m��p��TxG�~���T`Z	|�y�,i�l�^r����m��6Q�ZRS�S����c[��΁�'��;1��P�sj��"�RIs�v�x���X�5�z6�Bx�������:)|�ʎ�����ydp2��x D��n\�B�ﶍ	~Ү���5 ���6k�ƫ�o�6�K��0��) {������=l��	a�Jg �)n���)��kL�4�
�~�y��d#Ny��Ѹ ���\�e6��k���xC����l^kQ��~h�ꮟ�p����i�w�yGL�L�7Zj���^��cg[Ň�6�(KK��&[���l���U��>�qz��[�,1�#k���b�9��7k���"��-q�Z�.��m5���I���p)m���pA/���$_ž�O�v�ɡ<�*�60� q�T��ؖMF?��Ft6_��P��I�����O9�yo/�G�m��������Z�����*,cSS��Ϛ</תޠci��Y���?+�q*��z�7���{@������z�*Ԧ�<Z%�*b�V�4���Bj�#tnu!��I��맣_���ķ���o
n�O�9�uh���r'6��<����t��h���4��7RI~e�%V�i�QE�����B��˵9����ɇ���Ţ���k�S�x��gV}��L�hTvXԭ˙���������	��҆�U���O����w���(���g���T�]t��3�c��vs�x�m�!<���o kk�y�C�+�#�R�Ab$n����u��	�ꄅ��'Le����"ߏ?��0:�|te�[��$�E� �Z��e�9(y)щ�����a���FX�� h�  ��e�<^��k��y�#�R7"���er�"<��i@�<�W��	{�-!mk<��I�w�g7]���� b?�(����[��r�Z5I�bHY:� ��Ð�7�>����O�w��L���z�����[1�t�]�ٞ�	8_g�K�d_��=JJ��bbF��4"6��(��5�X���p3	^_�	�+Sn,ؚQ�]�>]1+��0c�X&�����V�ݳ��k��;�dF�Nϫap�.�� ���t�5	<!N��A������=r�����M��mR��U��T�}����b�93����N�����A�N�����V��}6 ��Y�}�Z�IA<!�� �B�w�������B�w貄%�a3�o'+��;[��ϲ<D� x<���]>y�(�]��y-�"���M`��e���s�y���ήp�	B���?�W~�zޑGZ��}>�ke�tɼ��T]�}�[���!{͇�F^H�m��p�#/��m� �Ѻa�U�|�N N��W@��H��a�`��*���S�S��;�C!�6�H���WZZojFOLM��ר���[�Bc��]�to�nG���@H��E���ߵP,��1�.[��$�sQ�)��FT ���#�]��6]N]m1���� 1ČH�I���qUԻv��َ��ehV&}��,�2ו���ɻ,�U)�Բ�d�6��پ�AK�-#2���0�w����>��t99��:LYgI�i�\��ώ6�_����+��bn�妢��O3f.�VA���9�ˎK4v�
~�b\�2�U���^#n
�R�%��b+����)���M���xY,�iz���w?�C�â�x��
���fSřz��H2�����_Px��Ti�`��K�0蛜�C�*���ϑ�/������y���3>V�L��~�!�%CE���3'���뵰fEbPQ<^� k����}{���G��Fd@�o� RA�.�p�'��X@:�{
�f� ��
*�������fn�i�J�;ˎ�Z�$W�,	m%�la@D1��΂���&˒�uv�B�e�&ݳ�@���R	���Yҝ�'�?�ݜ�0�5�m�N�+�S���h�	�
$�Z����>�	����+ψυ�}�&9
��˕�~9{��!�M(�Jƫ�P8Z�;X��M0I�/@�O���A�"!FV��D�̍�3<�����)�B9�U2��}�6�|�~y]a��t	k
��j7E���+��x�ܰxtg?Gś�����������[�i9}۬<beeu�8��Ց8_W=��u���̐וW?D9��>fx�>k$�� ������G�"k�"1��K!�����F�����^ǩU���s,� 9��E�A&�Y�Y%�,�+���޹���܀m3�J�HqW�K�J9
�}
)GZ��Q�U7E�r��w]�[e�߇��i�'2V	?��Bм�֕���D���X9�+=��L��~˥sdU��8�s�ȥ�"�tԯ��-������P����n>u�����E�i'�h�k0N]���M��Ђ�\�����/GA&Xșe���>z�Ժ��k�Htß8=*K�� �����C�*f)������&�f1ϫJ�A�`� `���͵c/_u��c�T�eg�\��-�T�\�^���c��vT��d���W�7m��;9���g��"�D.�����03�1R�#��C��|�1-
��W~~�<���צ�h��v	����#G��{�*����t"Fⱳ�wB� ����!25�N�"(p9cYj��i�_ �Q?�c4o+z殥Ծ�.bK�|�����ѕU�,2U���/���� ��������ݥ�1�F��G��k�ΗF4C��p6h�s�I��M��XM���S��b�K����wқ�x�����8x���ћ������.$'S�B���M�k63�?(�z�6q��>ވ��V�)+st��N�c+V������L^��ŭ���_��)'lu��t�R=����!��|V��#Z���������͘����ۭڔ���f�m�$,ۺȰ�"ޭ�QI�jG��x��*,O�������7`�LyǊ�;���h��g�@�w���o2�������z��0=����L��Ug$܁�L��l�)���hT��Q¹����4����{_�� z�����H�#N��~u��m$��{����^8/� ��?%��asc���u���H�g��T�tx,��5�3��d���B/ySˣ�p>�d[�Q�*;+��
�fGC���ϸ�ZH�5?�/�/E���wqsyDyT��-k����z|�@���#��5����g���At���,�\{����d��B��_(q�M��e`�6��1C���qz�!e�c�C�I���������^��`Ox+�G�6gw/�pj������)Ö��̒������x���ʺֱz΀�F�+��i��b~���N[|�v"!�䋨�&w>�����/��z�PR��=����OZ���f8�]�D�2����"�ݎ����a������7W@�G�oȺ�+҉rR��N�D&��x����d
� ��v(󆫗[�j��B�v�z�[�<��*�ի1Ȝ�ԳR��x;�+z4�ݙi\ǁ�VJ-zԐ��MM��<\)�dda��*��~T%�_�Na�_�ό���T�i�x
w��/:wwN�g�9cp�hz��#16�'�o��hg�����7���9��2�����2RC����$����`1�c��pa�����P�.��6�$U+�@���r� �\hF�?�=�� �Uoh��E��2�8���@���W����TifY$V�؂�J���Z�6��-�8��,2�n��% .],����G#��t�@�5�"+��վ�`��{eÕvm�a��7�*G�	��~L����|�R�y�7��N���������T�Yp��;��ue=q�	�&P؇��-���{�R�4�J��5Zp5Wպ��tq�+��K�(Ə�L2

�bw���ڡ	�2����h�l�W�A+���i�X���&��Vp��Ã�/���ȼ=D��Z��Z�7�0�GjAkfMo5��OG�M�c���<��:r^��������tg��2��&�cץ�-#i�=谻�������sH���,�Ϛ���"�-͸�l�֜)M�,]��Yg"�[rS��g��t~O2 �����ũ��Zo3��Љ�C�a�c*�'���ܟ�+[��[]�r��#��|�,`ņ�(��ρ��eu�Ț���V3�Ҩ��>��<��K�����������ҍ�j|l���!�%�nGwdhL��M�ef<"ǑU*��=�� �O��3�0]i$!@��
����W�X"D���TQ8�jtCL����Th�F��!���A����^�����d��5Kh���I�x����J� ��#�r���O�Qnj�չ�:�t������L�ޟ����ʰ�.yu�4�b�V���C�c	�0	��I�W��'"��������Dn��>ڢ�˷a��q_Z���Ul_=�y��w�=���lg�k ����o���(yL���[E�W\�C!�cu����-Ю�u�w�r�g5��1��gmCn#��9��m�yW���g�����M�]����=�{��``�U�Z��-~�?$a�� 0��p������R{����LU��Yw����G��l^�����G$�݊�3�o�Y���ˉ���z���c00kd��ɾ����K4�U��r9�.]v��h�u�����Pyv
p��tAIz?��u��!q�P����8�K��h�ԇ����-�7��Q� $�ۦ���[�r�S��K�����Vr��4V���{�5�2�/Ɲ+�žhy;�]�m�Ņ��|�^B�o>�N�i�[^���T2��$Y-���a �y����O�s��x�X>�U��ĩ�_8�{�)�:K<+;�Z�JW(� gi���?�? %�֏{�$��F�~��2fx���Hh�a��5�K:E�&kn/�8Z{����D
c�H�x��`��
k��:H��L�rצE @鋏���H`%~K^$�J�J=]������@j��1��[��u��RΣ�uZ��k�F���Y5hd<:=@�R�d!˱�%��W��{�x�p�F�!���b��n�a�\t�~T��٣9�|­��;�%3�-9Z�t�`�����#�i����l
�������ի��[m���_L��L ��5�Rͫ/+��~�^�ЪH��
;^� ^���RV���+f�����l�׃�q�YD4$h� �F\�R��"�I'������&�L,�[w�Y��	����V���Y�J�p%��4�v}�0C�n1�H֛r|X�$w��u����-x#=�)�i�FK�� X��M��8�K��;��eâ6E�Ɨ9;�V��&uG�e?�21�����`�/K�@D.��2�!������|��XL"�H��	����F!�d�tB�TU����������-�W�QOh��x���'h� ��1����� �ӂ��|��Te�L�
7�ͨ���_�D:��v{�Ԝ�v!���w�d�e���]�0 ��J�u���Q�:%u�(�CƟ����D���]��B&.�_S=Ld}vK}���$mT�o���� \������2�`JK�]U�D�L��-�3����v�ϸ�I�#���1���wR���>&���zI��0�T����g��R����ֳͺq��^�˵���x\�IDֱ�n	 �7)O�	k�}Zҁ�0����)z�\9j��|�$%�&b^��~�B����M��@;�B�=ON�թ�N|�À���V<ᒿi�"��~~��i�+'����ť.�%�� B���}~ ��Ɂ�{�4�E��O��
9}"js9�δ���]5�H�k1��s9����
�����������m�@bf_OK�2-��A(1r<��T�����%�a��!�o�~`�����̯{$wP� +�z��{̛;��o�����N��dӅ�얫z�'}����ή��t�Γ�`�U�����P!'#�=
�H_�"�֩�,T�n�0�g8���̢_��x)��ͨ�֬a��N�De5+ȼ�SO1����f)���SŔ	q*��@���3�Lr�Ծ�C�O���yg19�pm��2���9�a,U��8�G~�޿��r] i��4�x��^۟	s�J��*���X>#S�|A0E��"ߦ�=d�u/iU=Gq�K�L!U��`.4��XQ���q�a�8����X/!�F|pˊ�@~՛J�K��w&��Q�]4d�m�*9gx�p���$���)#
ԥ��aʐi�Fܡ�!��݀<���(�6l�Q��2J߅�&ӓ����	J>\<�5��mEă�]n���U[�+�rP,��u%#�n�Y.S�����,�'�V�1p��d�D�鮣H�E�/�y�!5��]a�4�ڑ.Q�PFq~�,����QK\6�I�9Ԋh��gb���󤝔bxk�R�ꑰ�ǏM���LJ�/]�'�|�v�B{o~�(=rq�J{����	���yV`�O��j��!]��O$(�k���/���������c�l4�v~&P
#�4yX������]���)7L�eWY�͇�x����O�-HD�"�����Z�}����Q:�`l�keS������������8"$��8��[`�1v��g�&�y@��-�3yf��q�K����-����<���+���Tuݿ"Ԉ�cKf9,��iͶ�1e��-]�_�٧��0K��c"y㙄Y2�aAؐ��	���#F.�߼��y�5]��&>Y�	��/R9?ޖj72I*J�`���Je<���t��e�1��Q̊��к�x������|xuئ3(��_���Q���\ʊ3/�C�Do`�V4�o�u���F���ʷ�D[����*�dt�
!�dfv`Ҏ�I���X�����ޕ^ ��� �'nn[�����NF�t},�MZ]�%�-
��+����`#�r_+��.u�UJ�~g�J��IQ��d�ϣ�򌣎���[h��VH�=�-8E�-Y�.c)ڰ�0j��Zh-�L;�8��j�� w��F.d��8�Ss��q�d%A/�Pʏ���l�Z4
�(�*�c��i�AaI�I �==�[j�G6T���K�91Bb�^u*��n���4���+ְ����C�y��k���w��l������I��8���Y�^/����E$�x��D�HT�T�f<�졄������C_�S���t8r��H���T)�9����~���$���c�뜩��i�e>L"�Il�S�P�O߸#f[����_�����.�� ���a�������������<�,�jY��,2'�� j��I�;C(ڎKDf�-�B����ߨ�������'�:8��GkX��>���O1�����{ӱ�B��d�H3տK��_.�M�K���M\�O�G���ΐ�s�?ěo�QX՘W>.[��g�=�;��I��o}#5�O-F�2��	�KC�"��OA�a��g��&�赿Q����tM��e�o�&�ޘ/�ji�Z�c7�:��[L��	-���T\�ڛ�ѕ��m1:�����c�>2�\��r_K�^����[-�δ����Qy�M�|eYx�AF�ܳ���uY~�r���t5��_h;0�g��";Y	$�݅��x���	ky�ZM��	fG����؊y�b��x<>���I�����۔��I�/�L�H��yi�F�gQ�����-IV����+l�U������՚������>�k{?��������!i�����*O�8�p�&��fdUO<+uү���V�P���mݞ#����h����6ba��Yk��>�vV�sth,Ͻʍǫ�o��i��+M�GR�&I�v;b rȤ��*&���4�.䔇�I�^��P�+�{�g�C�bf�w���'W���m4���^I�ZŰ�����\I�"?��7����!m=����~8S�#���L��������f��w�������)`%z�O��ַ��\`�	��[V�i����D�7u�roKj�"�\�~�>'a�z	��&�^�n�-�g����1w ���Ь7{(Na3������klI��x�
QJL4��iA�Hw\[���M����)�u�x�ƕ�~��*�gެ�NM�08~L�˗h����l��!v?Uk�b�@�kL
�}��G[b sLe�l���3[���K�l����dB���5`?�S�L���7jC���k�Z�*���,S��.�G�:�Z�����-���!���Q̇#��_)^$���G�S�l�wi����q�e���	�'Y�P�����f�d6%ÖUR�)~Qe��
 �.U�&D0Ĕn����|/��g�aͤs�SCaaϬx��-�PY �!�aJD��p=��ט��a8�"��v�8]�vX�4L�1#O)��Ţέ#S�#���G)��h�a���g_�0�W��[�(êV�#P	����d�W��ے�m��o���Mg�k%��BK^�$j-5(f�6�m�~)���~����P�t^ip��u�=i�p���H���v�T��Z���T`ڨ[��6
}C]�B�PZ���ŷc��}ѭ����ջ�np�~?�d�Q݄��rd'�4�GT��	��O��*��k�c0�4�G� �-��E_*<���-������e���P9>�m�ef�&���ZY7��m�?����&Y&����͋�P1ľ�q|j 3H}�<e#b�7��v�|�~���I�������D��s�츴*\���P�ә�#In3f�H�]����c�zb���xz34��l�,��W�����K�lkB�q���o����~.1�Z�Pڳ�O��^c�+%mE�0�Sm����c$�>���c҇2Q�����<��T�S�bDR����a�6kd
��w�G����<�����b�W����)��,��˖T�����H����E�	}F-�!O���b&MƁY�������ɇ�Q���=���uO(MĎ���'���I�����$��V@.�����RB�6��s+ҕ6�袁�,R�@�p�4�(����Xo������C���{�]?�;̲�)��f{���h�:��L�c�W�3n�Ӫ���L�r������ժ�R�g����4�8�4J�+W_(���Ni>4f���l��~��f�^�9�a`�c�q�!��.f���(���Iƈ�5O9����~����DsU]�r]]Re����%=H>+� �#��+���3�;kN>(Ω/4�e��V9h�d8J)W��ǆ �F:����,v�LQA8%���@��Ȥ {�R�'a��ƿ����:�s/�Y�!�N�"�G�{� !���wM���Xu�۔ }$�λm��y�Xk���#n\�'ۖ�� ^��5�EY���d��������`�2����H��`�RHj��>�����4�pZΟá���nB_����ɋ���nM�h�DVf��|����[�_20�#u;4���]B�?��D|b��x��H�Bg'�s�ɤ�G* .3��M+dA='�g�d�-t�Smfgu{����_]bd�R�"dk`p[��Ɉ�y�Ë�ޘ���-�-�cU��@9��;��d���܎����Z���{�A�1������]��E[t���(���o[��{p�=B�L<�G�N�Eé%�
�����V�i+���;��nj���o�O�J���f��EC�[�&^��a۩��i�����=�,zi�,e��;ٸ�L6�B���rv�%Pv,�"�v��6[��ha0���?��E������Yļ�sY�vF\*��A@�����C�(_J]�"
�~�}�6Z����ފ鋼�:U��y�Ee�i������ ��s��s��sq��j��gM��"��_���otO�*2I=aU,<��őJv���5�oQߡ���L�1v�Zs�F4����%����\E*��phVF�:�K|�hɪ}{��1�mZ���t�3��a�Y`)�V��8�6��t]1[�Iچ���(���&��]��X���D2T̷�LK�c�ހ篭u��Y��W�-�і���5p`�G�9אַ��=gcv�S�_FI��sp6���ڤa~�A{�OԽQ8�!��H����h~f�F��[���P���kM�-�"�'$e#V:��{�6������8�� �}z��C��AB�[F/QJW���Uo�I�������r(����:�� 
z��u������ڿ6���������zU��۶'����``�h��t9�D�
q��e7htaȲ��կk0�X�(R1OA��b�����w�ˠ�6i^@%�ݰ���t*�D?5��/.%��~/�β�K�K���^��Y�]����ԯ� >S�ux/������ϔ��� 5һ�WD������߹����t��oIu�J�OYɣF����(͙~0�ھ�)��R%�VY������e��ЁQYZ�@��&�&v���$�5�]���jwv'L��e�t:��/�(յ5a���I����A�[�ߖ�ў>��gcQ�)A�
�rz�e7�*��L
_Pr�!��'Q�1U�{D�75��k���r�[���{��+��\7��$6.��E�/F�!��o����`����z����#�����$�
�ܧ���Ex#�,�����~'M3�~��6.CwЙr�+�W�gZ�ШK�_�����IlC�H].avq�(�63�]���r����h�/�n����9��`:�/`@gI:�^s�`R���w�����R-�@ktGk�3b����'d�Rc&'Y9v��@�<Zu���,�V�K����<�< J��<&%Hx�ɡ ���
%zS��j����dI��x�	 #5yN��7Y�m/(wx)㫿�0��Dr.�≚&�@�`�)b���֓�m����x=�
tX[D��F��^0�^o%��xi��������?���`8Q1���25t)R��D�<���4�js���#p&{���e�j2�0u����(w�wɊ�����Zl*��}M�>kN0M��U��/��'�|��b��2eM�>Yjbo=�_D�f�d��Oe �BF�tBF�@r�t|��#�7��M
o�)7����r��p���-^!�����Pϊ4�ѿgM	�)����1�����0�μ@����;�p�����e��n`�|��.�(v�@������P?���>BRZ�L ��m2�fK�w}���m [!���UPZ$�ү0(vk���_�IK��X^�m�T�����eW��ד"�R����$|�Q��U�4XW�� �{T9n�Dao[�����ӂ�)<􎬅��Cj��|д����AE�ʏ���i��U�<�TPt��/s�]~b�ci�r&�6Cz����F�݋�M��N��p��lw�)�T7�n�*��q�+:-l���U��+�J񌴫����K�JCI?�~)���%�|v�H5m�����>�Ŝ��cTm��8fo�{|?��nziIg��D��2%��N�@&��Xƞ�iN�mAu���6�z���{�~�X{�w�x�x�X��:��:kF�; �q��X#H�{��#�T±F�)z:d�*�9��52Z�.1�?�5f�U�_f�ʑp�ެɑ\(Y>M��&ǜ��qJ-�XV������zJj�/�q��O�l^���Z�H�2�����^B3��M9:�p�,-�v����2���*����e̝���Ȟa��b|u��#�)ճ�S!����}� t�V�����x�@MTS��	�R2=��]�]ί��Q0#˟��A$L���7�e{s>@zVó����q&ex
~���)K���5
���Z�o�&�u���x2)Ocٯ��pI���e��1��~�7�?���!�)%Jz���ߺ��X��%��3�B�vp�e߯�'�P�TZ�|�YO/�(65KT���0?y`�q�O*	uj����|��mN_�|+��s���N��O�2R�B��S��;~���̷<��r߶5h�!����x ྆yc
�����:��5^�W������v��}�{�e�����b�ˍ����ƌ�=ai���S+.. ��]�xnI:+J\����� ���r�3���UA�V9��o��@&&�\��<�o9���&M�惮��}���w�d4�۟����ŞN��l�p]Ξ�`�@XOղ.�φJ���"K�ǍJ���>cJ��N�K��Y�ә������|c4A>?�N��׍��ա����ڕ3�Q����N��D
s��ct�g�k�7��r�L�f�N����haV�~�^�������y�[O�|iT�
6
����I
�}f�P_���K�F�W;w�Jc�O���X�_3Zul3��ԗ����*�u��a&y��w�г�Tf�z!���4���� ��x�ۨ{�3k�n.�f4;D���z÷�O�c>y2YH����Aݡ��0�694Ʉ�;�^�s�ǭ^~�]��vc�H1�
����C�[��a�|�J�L�=��9X:q盽VW�V�Ϥ���-3���B>\Cm�?x<���Ηg�<;D�1��|��qvN�H���8�u@l?1�l{h�60��#��򍍥���v�3\攳mTs�'#T�a���<���n��^�����k��{u�&v�J�wvR�/�}����g}�����_!:9��n�D<7�>���!���@xx��j�[X�������i�� oԸ��:��h�a��o��e��y���ei�+�:�����i� �f����<�>i)�k 	SK���[O�-�e�6��Q����C7��+�C�k��جZfNH*e�2���Å�؏�k���	�
1�
/P2��\z�{2�3Ӽ��7�Wc>W��"�����94�=�4����AK�,4����I���&�lV�C~�[$2��평(�$K�֣m����V\���2M���b}�џ�g�J��v����+\ٚ�H��88��T��ʚ�����'m>��$�H~Y[6�Z�Hވi�Wh�(���º�w��4�2�2#96XC�>���R?C���G�4T�I�df��_�$�'��P�nQ{�aT��<�%��|�?�aq�����ױ�$� ��ߛ{KG��o���'M�?�r���/9[�,M���g�+���sK�����><�Y��i��p٦"ݢ�&D�{S�QZ�Ն�LsM�ް/+	i���R6���dk�G��.<?\���[��ſ��:/zb��0w�}.F��4.f��ӆ�dq�YĎ�)O���C�L�HF��TE�zLb�)-Y@�s�m��FPv��ɡ[7/8�w�x���s��d"6�"�y�2�?��"�<�BW}���2�K;m��Pg����.CA��<O�A��j�bx���i�/���f��i�2��TB�J{�gjt=��`s7g�e�-�_ ��i���a,/��	����;McZQi����"]e��"�������o�8�v �-��h���Ň>ēK-`f\����$8i�u�zsU/��T��cS�%��m8��O��,����]�x�R	���B�
��zJ�yv���uF�����'�YA��mSA��v%��q��3�)�X��\|���J� w�������:���J\Z3T�m��_�gt�2�Ϫ�+9A�G��ɚF�_�U���()�Us�^��-��
�%w�+��ޒ�?.΂)h��� ��Bp��'���6��!H�������{p\���S���?aKu��{u?Y�Zuj�땬Tv�+;��G��~��3�2H�U��=�=���"`?G����8r̰[-��'�	�_��>��q��=b�� ��0H�&>���*8�S�籤G:��:��t�+�癔�O�:�퉂��x=�3�s�Z��K	cM;o��������K/_�$9+�r3���6.֑Dkֶឫ��a�:|{Ī��贜�^j_��8�5��ѯb����R���.�a���8Wc# C�,f��E�~����߮x�.xl˒ܱ�D.B*�^ݤ|��$���o�g��Z!���� Q�y���
�u�
X��y{C����XF��B�k�R�)W��g�>*�$V�!Ӑ�+���"5)ٰi�\�bG���`z���|�����׵��l��r��x���6�Z)��W`F5����D>[d�:w2��Y,�<G��,1�<��(����݌���>������KjU!b�X�SL6�P�~2R�/H�É,Uo��۴�b�'�녞�i���Luxidf'ld�U���()�=L��4PI	7���6\Y���:��ױƛ)�c����[�����������\��9w�|"k�9`l�K�:Ο��k��O^�!yo�-A�O��������O��r+$B�M�8HY��>��,]��3�#A���]�5z)Hu1��Hz5���b�Pͩ6�6_�_����oyۄ�W��=m���S�_�h!��z�lQ�^ !*�v��g������Wt�%�[�Z���q�p<|�ت�8�M4�s�T$R�u\j`˃�\m���>w�8��Ϡ���t�6Eg���̠ݬG?||NdW�j�D���RJ��vG��M����u�����X9�������=9������9��ǫb[�(�437���(����n�Ǎ �&�oG
s���5���Y�Gi!�\�PC�P1���!���9X���kS�\�V���^p�x^�O�Ზ*�A��O���f݂�4��L���ʾ�el��mv?�<������l�Ԝ����Ƙ�ѵ�(���gH�_~D[ʿ��&n0������ݱ^��c�G�@c��»�Ёm!f������]���>{��K�G!v�����BuM�X���W��-���m�*��Ʈ/f
�O/>�n��,Rc[�'���7������w`�;U�[�a��=ͻ���Y�a�/^��g �Y�V+�b[�r�2F��rxO'c�J EH�����@*F�8��.�`QX`�\�XLG ���8Bz�Go�}�,OU�1���DP�BnA��I�`d�Q�����MvGD��z\� �r4����K�nPQ�������C����y�q�>;P�H���P���ϑU�XE�7~�f�lTp��EH�^�mh�+а_��Y I4����s>�N7�c���%/P����7�$E-1��1�w��`���H�p�<sιW2d��X����8_��p:ڸl�n��%�&���w�
Z�~�Z��H�!�ц�b�k1�՞ܕN3�����,�	>����5��
x-TM��?�		�([U��U~��һ�VabYG�Ref301������u�I�ۃ����������Ϋm;�R��/ת�d�н"�����煱���;6��k�8��3*�9�fr��k��j�X������i�qL1$\+SY��D����"�Ū([e�̂~��F�ft���0�o_����Yn_F��1�Dɓ<��߇be5����F�����Qm��	XRV�����w98�-@��2�]'zйwŢ��M��1�27��~8�5���`�˸�|�s��n����c�q?���gu]�O����2.�d��9D�������E��l�b
�}cνӵ�;�����i�G�ӱ�ɚsOw|��D��Բfk�c���ch?���tB�9v���� g�S 2��*6#�	Ë�+�|����UC�?�McS3_c��7`xi�8�i�zP/hw���d�F tr~*�WE�7�PdWY-t��h�߇c 7U�_D�����p8�A�1�p\���7�[�3�ԅ}y̥�"�v,��Y��M�������҅�Ǖ�@��293Jr��Qa�����L
��-kNɘg����1�uf>�+�� �J��s�@�0��q��t�a�oo����h���T��to����1�r9W��>�9���w��iH��4[yӦ�c&l��
�oP��AfC_YD�
�h�KKىq�#�d������i)o���]ͱl����:�+��sp%��1lׄu����˅��s҄j�V\��_͙3�:z����!ԟg]o�f��%`RV�&�U�m]�ʌG�R���5ñ��%�T�[��������Q�I�B����>����O*�W�(��Z���7Y�׎xb\&��Q�L��S��5������8���w�੨�ݽg������=��aq�nh�U~NXU�C��)�����q�n���a~D������nr���t� �y4��wi���A�(��z��I�ɖ�6��QQvv�	��J,�������:W:���0�q06�_+��{�@B�<�K	�FFp�~�F�〫��f����_��l�?!2�@�]lۣ�[�hT ��`X$�w�c2��/�E>r����̳���@9��e�Fد�O�t�y������mش�*	E���`x��j����	����e4y{}�Q ��fkt���ᙬ��?�-|�C�p�ޡ��r��.Sz&bBA��1w�S�,���}��B͋fx�ٴ�>��i>�G�M�7�_�J�(7`�P��,�I��EO�[Tkt��y�~d��F^�����^חb��˚�DS�����iw2�a�c�<��Y��� ����r��U�_Bސ����y�����F-]�������a}�䂙`q<�%��TN;���L�#�A*/�c�J^]W��@�?�d `�O��Ƶ�˶^:m$�Λ0?�^B�/�i���gu"v�2!���@u6ms
��Y���2nK�P�ά���e�?+�N߄��ٕ����}P	�1L������� ��KЦ�4tQٙ�����~���`��~�og�5i�ҩ��8R5+��XF��caـZ[i��QŦh׀��Z��l;��U�(�2\��？E,4@�oZ����v�O��̎��vElIw�K9�Lk�o`�H�w0�ϟ?�̙�'�'�k0~}�����`H�mM�f7���5�1�{�eq8�������}38%�(�r�/	|r�b���2�Wu��?)��}8�@�[��Lq�e�9 2�*��s���r�#粈i� �I�)��$>=�ׄ��Y�}�߅�u.ĵ�\ƷL2���κo�I�|O	-,����L�e���1S��05lt�́�=1r���߀�PkM�l$Z��F�E5#�	ܚ�̊0b�$���G����^��!ZzÔWX�&�!�G]�N�c{$�����{-p��U���}ڱ��xz
�ݗE�x:<��r��Ǻ�wF����a���o;�2��{c�g���k��v�q�ū$�@1�"�\��=ɛ,�Ѯ��A��>~�Ρ߆����8�͂E����i��̱uf������>GX�gi����eh�)����ـ�mo|��-eB- ��h����'J��s�Y��?jvl�e V�Y�2ix��&,�[��5L����PG�@P���{wk�w=�PK�F�6z)8Ԍ�n��N��x��>�}i""�i��;�A���c�� m����Vh��C������&��h������:Y%����
�VU�Q1aZ�ϩV\�#�����8�Z��ߤ��o�q�q~C9�lba�P\&k�$gk�W,Zwߐ<2Ϥ�q!_��>��ݰ%�H����6jL�f(�^O���N:���p|�h����˚C���І���p����C��xPJ���Y'�2�	�h�X�f�D��L��6m�<�%�P��%Tt�-%xZ �h�db���l�-�':������d��Yx�ZW�w��AlxH����p�����)k�4v�j����eK#-1_�z&v5��� �����u]�ˮSyCŧ1~%^>�W���ױ_���װ�;z�0e�Ĵ�O�g�ݯG(����߭r�E�?�oa�oda)��f*�ֱ�E�nU���Dَ�M	S3ו%?��]�b�%?L+���G���QQ������z�<_����wz�Z�7�Q�І�n��ܡ�1W� @���9�����L
�45���������� i�ⵙ�$f%-�`r[E�̚mɜ�;���3��c��	����͹(Ʀ�S�1�k��f���+'o�':=w���R� �Q�~o����5NR*�
T�3&͢+������2Ź��F�gm
Y�tn}8Nә�ّ���<�C��ɢJTl�_Dz[$�:��]�H���:τ�V$��w��g�ܳ���Jyؽ}���:����锥���i�Y@����B�L��g(����C	�&�WiY���u�#�i���s��K^@CCܾr���A��~��R�QdP�j��;����aƳ�r:�Qe�|��%&c����ǈ|��s�5z5����y"���wr�_F�SD]k�j��ũ�e�|��輐3�X! �7%�>���aK�గ�-9q��_���J�>�h��<a��d�m��/v,���Ili����l~��3͗Y3g�U~K��{~��`�On��Ͽ�.��}+���5�u�NL��_��"N{\���ڄ���p��5�?����duUАťMY �f;jN�L܋&�V��M*tW�_ee��wmF��s�a�c�a(�i���S�E=��U"UHڑ���euT3@�>ֻ:MuԆ6B'��k���W���
�k�� ��~h��
�[���&}9�����V!0�+R� 5��"#��$��@�nT�Œ����
�'���z=P�I}P��d�Ҁ+�ȍ.�Fq��V�a�}28|�P�a���SoL�u)�S�P\"e�Ղ��tJ��)'�B<�)�����[6�� �H��kv0�/f�ll̍�xN�x1䱣*-5�"ڐ!���uaZ�;ks���>�~106>1*�V�e^D�5�~�Ȩ�ԋ�^�����(�ŀ�=耘�B��`}-6�FX�k:���:E�Fdw\WDNLP6��	��8��^ @'�灐�<��������4S61 u�����m����+f�,X1b*U��H���] ��U�5����3���WTh���Pn���a ��R��A@���m�=m����8��g�|W�rg�UFS���0J�MeB�D��nq��J���ic�I��|�
Y6��~��{�*Vα�U1�����\a�4?��CH�C۾���-̯���g|��M�36�ݾ[WXW����'X�\o�
��7d�dJ�����a�ҧO�g)��VV'��F�'<Z�Á��&�e�� ჿm�7��r�\��-vs��¸���r.}�2Q�t~e�%���D�1�����D�xc�$o�@#ұA��6��i�0|�E��a�4k���I#�N����f"��%����W���I(�O3�r8��� [���u�@��'�J!�,+� u��p(n����>/y��-rau�oȊLc��Qb������K�<\���MWsU�a"Ȑ���t� �b[�|0]~ɔP��88Z3T�S���vY�\	X��ZUkOݠ���.؎����\�4*G�P#��Lq��V�+��*��������ȇ�v��U�� g�I��'_G��2&Dm�bVp�&�A$��j��e�m�2}ʋT(r��7	1J�ܺ~qm~J��&��	^�:6�;׷:�LR�b27��P]� OX��s�ށ�&��X�Eg4K;m�򿘜~����>D�A���W���$�vmW:+.�>h��P]	�~MO��1�~ݕ�0�q���\ҽ������"(���ߍ�L'��|�=�;�XG�P�&��%��X��,�����n�d��wq�|9[x7p�]��~���n�+�q��n��ñ���S�-�ׇ�T�?��jk�q]�%L��[m�d�vV�ҜzK�b&N��ţ�TZ���\��ѢЮ!�C�Mа��$g��~��N�\�^�H#�ܟ����O�$�NDR��+�i�O?�q%Q�����W����T1���ɚF��>��"O�u� 7���~�=��?n٭ƈ�� ����,��;@����� ��:F�y�O����z��j���	 a�*��F|�j���-o�G���n�a�R��fr�XJ�J��o$�����Ө�<���>6^0,�*xP��g�#��P�D��,h�!N�ۦG�6|r��?�a4%?�/�<N��,>{�댞`�#��0�A���o�Y�l�j1���"��������Cĉee@����:*@`�{X����b�*�B��U�b�q��V�Ԡ�'ǣ�>�ҙh2сV}�a�8I��v$�S��GH��4G#�j�mQ5�j���*쥲�w�ܖ�����E����=��ousI�A
Y4��hq�n�en��?n�K(�_@��u��-����h���C�խ��4zXj�:J�����g5����p���w��XL���������i�񲢗��7�`���7i�ykd2@N�Cs��@���zpm f@�6��Z�%�s��	7�Su5��ylND��{y��ܴ�Z���*C�=a�h 2���f��X�z��:�N�"��t��ͭ�F�-ݶe�T��af��Q����R�a=�! l��y�����/���&�ӱ��ޯ�+=�TON`NgxW8hV~�|��ˁ���nb��3^��?�P�uW��!����Ձ�1($6�\�Wc�9���~K��32T<�ju��Τ(w���L��-v��@��ދS� @!5)JA�V)kV�鼼�+���kʧy����(����W(����a� l��S'��뷛��M�SMC�����!�͆��� כeh��ֆ�I񏳗�7��M�۔�:w{��-��T�^>hm'���>飛��S��I��sߥ$ ��:u�:7�1��	O�$�[H�-��L&r�GM<
T�R�,V����ڠ�bZBd�������RI��(m����]�����<!} ����v�H6f)����L�"���m��5����|��E�S+����hD�����M Z]f8�>1�̹�i96M�x�bc�!�c:�L�����0η:���|����}�� ���_6&k(��.fp;�R�r.%@��C`��n���L��x#mV�E�[����Rj�;�h��� ����>/E��E9F�.rK�nӃۺ'����A�B���dl� ��������p�>o1�%��"Ęy�o�n!*L����I�Z�> W�[C�SȰ���"g)<6�N��������B�w�y�i4\��3�Hʹv���Ԏe��ݟ�  `�ngD�@ k��EtC���DI鷋<�2�B��jd���g�r�y���[QݝD�/=�?��}x޷�^��s�W#��wKWS-sa�C�bOG/|�O�YD��5c��_Vo�K_^T���5̗Ĭk��@�P$F�}M�N$�<�By
K��2�ȓ�J�`��R������
�l�<��L_Ύ.�6"����.��4t�yݔlw��|Y~���Rдy���|`"����0�|Dr���?�2K�,)8j���5�$�vC�z<��`m��Bt�[���p������S��B��Ѣ	Cs��m�4/6U	���T �ET�2�V.#Խ���ʳ����u��O?�Z)L�^<�D�r���z����~
��� �vܾfV��c�':�]8�Q��O!���w!��Ԡ�h,�e�We����s/~;[�m`�0C�96Q�,��6a�7f��-q��UX��{��ؾy���(����5�Vf���gN+��O��]e�#��4�c���E���)	`���񇸪%~s���"�c:KZ�c����/H�;���2�uF��?��OXl�H'Js#��й"� 3�ry-�P������NI��<%��m��Me�����cKT�Ap�ݶ����+v�����PF����m��]m1~�����`�b�f�<Τ'f7���jӼ@7u(��鎢�5�h�ݧ�������0��mŉ�9����ή���^�k6�' ��g�u�F�F��;z�����C���̧��sZ���y��n?k�Q#���:�h)�:���2�"m��YL��oI��GW�J%��&�����zt��I����n	�rE����\&~ ���DQ{QZbOh>n� ����#PWb��Y����:Tѱl9�o��8M�[>�����"J�y��Յ�T�Dfn*��N������mZ@�d#Ď���*T���b��Mo�b����V�6=��l�X,�C*����N>���`�U��7���S��������,x�ԙ�(M9V׉�=a�!#�֜Q�P���e��g�bs	D�[��R������^���0�m=�=����]bJ�\��7�B7L�;ΤH��${ �x��`�~�!��<�ۺ�d%�'�a{dZ��@[ɆoiɪUֻښ���EGMa��	���["Ѱ���P<!�����F�x�?r�䭦�AR#�����%�4��)/�ʠl�0vY�bm	qLI��~��odW��{۸Mkw����?��p;!������b�Ф�.�v2oP���t��>���(dT��A1�?����8|#Fy�Ќ�U�Β���gW'�|W����/o����l;[��t��c|��O�C5m�2���+�A%BfǶ�y�J������#<I�J�sR
�Q�,���q�yk�W��r^?`P��߇�{���޻�����Q��mo����%�v��J.�wT�_}WJ�(���5wڠf�.�} �P>�J�r���*�L'���G��ɯĥ�m-��)�s{�:�����G��H�9��4�}��}��(l�\��%�D�5�%�l��\A\-2��g ���-q�[����@��;��R	'"��Z `SYQ�{:�{���x�ȥ�I5�����oPk�>��u�w&iΖrn5���r�965����aW"n��:j���J��φ$�)&��ʥ�N?!�Mkx8�[ w�̞��1����e��EL�.��A�G{Ӷ���r���S��*���E˦4c')?���KS���D^~�����t�Y���;Ȇt/���o�U�mx�r��G�Ĥm��-��U�G�����/���CNC5\�c����O���P���A��S�ک��q�T�u/����6�"�ꜘ��4�ȏ���7|�^:��g[[��j�x�ۚ����^l�^S��G��wЦ�������7�)��U���l�?�s�]	Yu1�k&(=o��=��V����:�%���ˮ=�BO힗p�p���-���c��b� � 2�ɮ�s��9�*n�3>���}�&�A)m�B��l���r7ESA3�Z����]��d[ɯ��m������ܟ-�q������0P�%,7��y��5F>?������6��%���B ��;���
j�30����ߦ��\��/s�����o�=���6@�yl��\���}pq���ƕ[PmX�2 ��P�. ?����i�o$Т`�I�qD܌��6��(�����Ȏ>�?����$�K+]9@�Z�߃R:ڰ�F�+So�A�ÌB�J�� V�8"����,��ϑ�K-^�+~3����R���M/����Ur�;C�ר��Q��Wĝ�'>�Ƨ����(I0�m� A&��25X��w���l_�cVC�zJ2���i�M<��w滙�JV-*����Mgp�	�0��W�4�S����v�u����F����ǿ;Ij�_̈�H��*�v���*�T2������,����c�`r�A'ASg3�\N4�H�݄�t��}�\j���_ջH��ew�1�}�U�Fj��L���_��힓�ޖ=�$J+ded��^y������\�Ƭi�+*�^�D�V٨%ύủ8�\Q��S�6?D&��=�Y)-�C�jx��#9��˙R6ȑ:&�Ʈ��p
�kDj�9|V��+ј�t�
�wfBY���JQ�y�e���t�'b�[�*��6�@v�J�Pv>�@(�|U���� �?���h��A���z=5�2�Q���� 9I�N��yZ�}�M���>��v�i}ʐ��uWȺ�����~"�Bj���W�������q�}�Y�����O	;A-�r�)|O҄tՕ�eQ�����������~"��q$����U��1���Y=���%�GĨ�9*М����(�����VHc��l�u����e��α_�1?�� �/f�`5�Bmd�c�_��b��k8o�wG�.�M�!�N�B�`�6!�P6�H��ֹP�wi&vN�2HZR��
�6�q��L��lk�&h��KI9w	��9O�?v�z?����Ԣp��Ӽ����>k����I�{���Gc=�8��ׂ-��lcee���G��)Wa�zן����Oɦ���I�e�Eq�J���V��d,�T;��VnBD.'x����ͥ�ҽ���P�j+���5_��'��s	�O�lB�y�A[�=Yc���>�o!z �3�x/�^�m֥����6P��9��LС.��i���A��]F{�G��H@����p�.��蕾�~��RK� Wzq���D�B4�휳5�i�*M�m �R�lH�o���(H�%H�2(��#)>�	��i��"��t�x�dk/\��� ��׺�V�cwyi�5Z	-`N�a=����ѭm��F��GYz�_Ʌ�"�+"+��3�bmJb�"9q�M���t�h��麟���<1�!�l�Y	���_��3��b�~l�]������65T��T��RȫQ�����{�$�Hｾ�銄��)?�T907���fq�o��⥋s���v22�k�)ba4[
�QΝ�a1�#c���>S�,�;�B�v'�3#�Kg���3�tCY(����U�d�X&���gK�T�
wS��_�t�Zβ�P�3���,�l0E���G���!S�j�Ϊ�3�V
�z���[L�/}ﲨ��of�Z|1�}\l��~�� �Ot�0���Wh�J=�mj7��v����%�Y�R`�h�-%�ӮknFdxr|�ByL�XG�l�����X���|%Q�=<�O�����0�xmT%␃�Xv`����Y��c�B�*4�-'����o�젼^L�;��y���ն=6�oE�0{B?�{���\v���ݵ�Y���4'�k��}���Z$*�9v�,�[ʃouph��b˾7��E����w]f|�4����\��X����p��k��s������mX� �#�E�S�f)�ϔ[b�Q�9����M�S>V"M�d��T�>���F ��B��c�ת�x�W4*����c����/Smp�h`a������\T���ᬠ���/���f]-���i$=�lP�̽V��Y��T8�~��u�ܧ��X/Q���|M#��>&L�%�����p��凐�=��lL`�צ�0l��#�%فe��b��%B��\OW���1��0!�t�M%6�(���E�dTL��/Y��)���3Z~,�S@�KYͽ�u���N3��& iAd�[���b}��00�X��)$�C(2��/2lE�*�F�,,��e�����n��K�nr����PX�O�+$z���'yt��K�h?�x+I�7�P�6�s�)��J�NSG	���*/K�i���%U��0�n[y�WS n��Z�� V�rM\6�1=}!X��>��ʨ��!c�3Pj�ف���J�;�0U�=��S�ʺ���bw^q'B��c��pf���f~��i���w$Qy {,�&¦%j���O�����G�ʑN>7��NOf�@0��H��'=�%�8���ѩ�$��8���]2���c�Q-T�M���y�|Y��GM������tf��� ��(���[��5pH�$�:Ya���I�#�h�9`��wl�U�m�L��S?��vo�GB���*�f�0-�8�� -�kJ.B����B#P�������!е:��r�im_֬�F�Q��1��=����0�R[L�xe�ʾ4j��ӊ ƀj�cY��-�r.�&���>h�;d�ߗ�5.ŝJd�^
�U��E��#K, GA�*31f�-�4�j*��>
ijz���
9o�R�^zK3_�}����S��ߠ��V�z���Y:=!�� �v*��M�Mڹ�X�,TR�ж\�&��V7Ԃ��_~5��mr���̐C����������i�Ƀ?�ˡ�t�$��@ӌ^
9� �r�7��Pv��cR֒	�ᚘ��B[�8��(c��̤�o���UQ
�-�fL���C�e���F���]:с��Yd��]sb�F���lQ{�u�֮��Fύ�rKv5�&�}�p$T����Y��O�`�aX}�i���%��ERtpE! ��L�R��Ϣ$_��X$nI4�k������p�<e�``By	&KWQ �
Ϥ-�^�^4����Sy�F,��ݴw�: ���}\���_I�@W�TjC�[[��w�Д����U����A�;�ת@dL\��n�l ��{�T��AD�x�~r�g��f�]9F��	0�!��:�B�]m'�'ټ��n���G�&���q(���	1|#��ߋ����3�|�5��3�D8�$8 OO�T����Y^���t�p���ޜ*�fO��I�߯NioԾ�|o2�u����/��ޙ��r)o�>h��?ji�2~��nC9"�g7����*���$(D7�@�����7�"�Z�&�d��#Ha,Z?��x��$�>EX�U��9�ý���pb��@"c#�������s�h�'�������5w��� 2>�z{ڍ$co�Ű����`�]r��͈; ���P_8j'�e짊��q�Pl��?Y��'��*�(��1mie$�o��J��:�3���Vx��!�&Lj;O?�ȭ�`��:�ȶ'=3%W-!;�S�:�߁���ծ���&����׻�iP*w9����!��>�ҹ���Q%q�i� ߃��_ECr��KI�8���뻋��	���`�������Q����e��Yp���bX�R3���x������^ ���:�Y(@��X�_^��66�����$�vOe�HA�_���Q�{���J��߾�E<q���f��M�YŒ��,Hfd��b!�{gŔ3�2|(��������`��|��`w��Y;:y=��l��A
��T;s�a� �L���hJ�*a*���ֽ.�u��I��;D��
E=�׬/��|]_�d9��n���[��h��Х�RX�8�R�Bo�'�#g�Q�Z�V�Ij��S�����aq2��._����:��X(��$Xp��I����������{�aÿM�p
�|�x��g��^����W�L�w?P�H�Į����n�]lwl;9Y��l����滛부S5����L���F�=�w��q�5Ps�_+�101�1�L%cV���6��8ݸ��\�:���R����nަ� nݯy�I���t�?����mo����5�5�r�S�o�y���	���5�
��ǣ'K'@��6��d�r��^�3��0ټ~�܌���#�v�l$+�����Z�tQ�Ύ��W�1�*���F��@L��~)C/q[�W����T�ʐh�ϓ&R<&ԏ�!D��K��(�l��	�VH��w�����y.���Jf��V-��{�۠�
�� �ϊ;�Y��ɀ���(�(-��ば����Y=����0������a����c��h����Q�&��-�=��x�vw-[ѻ47J�]��@a� �B�:�J�^ 2�e�k�{ �>�~��L�'ʂ�Z5#�Ŝ��,��vh�;�m�qmK����y��mW;�9�+ٗ�����&`�(�5�F����"��|�}��OҪ���	k�~��o2U[S��$�V��zPl?�����ҽO�#���|�T0T��i^�w5d��k,���G�%%DG��A��G�5���e�����;W��-�%����V�P���X�?g��s2�6Ѫ����y~ll�G��_*��fp���x���6Q�"pu�W�$�[J���;��r��ċ��㲿�'W�6~9����>r���h�Wa I{�`�,�
���K��D)|���D�C�?\��I�����^V>e"X�Q���<�����',h��,!x���G�����p��8ִ^I�7�����/���%r�zKsF��/Ɋ�Q-��@��xh�u�m�|�[=J{59��o���Ⱦ h :��.���{رUr8@D[�'��E�!������D�p�����.���&�.v{�ge����l�H�M�+ :<F�k����xW���O�m�*�
[qcG8�dHr�nS鴾�C�&�� q��I9����%�j�lGw�M���x�E������Ss�;ަ�=��d@nuC�N���o�-�ˀ�Ї�:��߽f�V[.*��6�d1��JBM�e;4�b��{%�=7��C�r�	,Wf��jM?%�$����_4�[�F."%ի���@�V{.4u߲����D�K�]Oߨ�j�^��,nk�/�m.9��a���t]?����{8o��*������$J�Mɪ/�Y,�Z%���˪])qҽE��w�I�Z�ƇrU��Uy������/�X3�EV�=�����+�$�x+�.I���8�t]탟[
�c���4)/�M�L�>�c�5sH����2_v�<�#�5��G0��Q�R�����r\�<��9s���^#)Y��Wr�l�F���ה-�v����#kf0��]_��=��q����o�&l�R�6���-�p9�rf�n�*�q�]��|G�Ã�m�6`D¡� ����~#f#d��3�U�Dt@�v_1�¢�j�+y���\Inq�F5�qA����A(f�����1-�XH�i�P��^�5(�)����0��������2U�o���m��:�o��0Mm�
����<��ue?R'�����%�(E��66a�uGl
6J5{<D+?H"O{b���W͋��?�09��O�q}{�$�t�79{�΢��
�:]�W//�À�v��I�B%9��nIJ�<�;;+�ʅ[�R��_��J��776(��_'t�c�"��޳3-\}uT̟BZ\�\u�'���ܤ�-����o�4&��ge���V�y�;��Y	�x��ۦ V=#�A����B�&�X��a=��5�W��5tY\K�a6g���j�q�
g�R�~��JN�� ����£��� z�6lw?��v;�
�!���g�m$������ Ԯ�*�豆ې�Ux]=�SC�
�\�HD�M�e5A�a��d٧u�>�l��Y��e�E��#h�����������'U�n����k#fm��*l���^s�1������ o7xx�7[Vb3y+VU�4HU���\���L֍��q"��J�8D�z_�<fI�N�}�����4�U�d(��1��W�2�EM���U<#���·J����Ab�R��;����Pm;��#�el�L/1č��e����� �`ޛ�����rH2�K���3W��&E:uf�@�� X��k�|�٦Ƽ�nۨt�Ų�b3��D�3r��"w��}#�4��4+�xa������t�ޜ4!FQ�Lg�Cu���B/k˛5N�i��7��d3{��kؿ�3������C�i��\��q=��7E4��_��Xj��Ԍ1�Fj�*�Ì�rc�ۡ�b�]��]�F�g�k��z�hO:˘�`�"�Z䍓��@_W��T�k޸�f�I)����UGZJ �}�Y���ߍo�7�s��d�BZ�#>��G��1��ŋ���Kn��W����yۃeOW�b��u^�����5x�D�Q^7����C��(���V�,��adK��ic�k��#8��
���x."�[bcf��e�e����u7
WYJ��;��×b�l~|��Jl�ؼ��wu���/st��!y�Z���oN�~�"�ZJ�S�Us��᫪�C�VB}|��<t}�.�'��!F�ɘ�V(�fi����)R�mr�">?M��4k�I ��!^������W�}�7����O^\[֞�_�7�O@e���DI	����ǘ�H��~����%��r��r�Z��?�o��9i�����׳�l��;���v�2(����x7ָ;$4��'�����M�<��qwMpk�=xp��;�Ss?�יzO�/�j��o�:g��9���%>7{��Y[���W��6��M���[��>"'��A:èC�X?�H���	�a��u-~��B(uh�%�8��Rܰ<�Z�X�����~%FV�t�M�*�щ0�z��:��횼D�d����M���Vy	7rd��j���kÅ&�SKj�P�����7�5Ȟl��vK�X��/�+?i����O0UE�c����kV�̬V� !�XG���@gX@ۑ�PV3�A�ք��nƂ�X�qM�F��Qv4�)|x�z�bw~P���]�֓�o�u�+5�0Q�v� ڦ˪��/B5"�Q����ڦ�r�6�+Ѕ��1��g��L�6�T�"��1*H����aTWU:`��%�Շ����3�����&[>�f<++pFb���DT�ȥ�hp�3SR �7Q�Gv`�����qg���A��)���F��ԯ�ۀǎ�V�p����f�L�4���ދ2��yZ��LXh���o�S��] �ߕC�dy�Œ�dVJV�Z�bү�\�v�0cM.�&^�\W����s>��칈]���He���:p"fh���+���x��c�J�	�O����ы�T��[�I`����u!Yu���}��M�d2%L	�Z2~�A�֘�)	Bp�x�r�� c՜pZ������|I<,��8�C���0%Z[̈��Cر�T���C�����Tҳ%��	����`;�V�խ萳X��-�5{�*P"Cx�r�_y�%j��3�B�e�.]�`�?�M��9\L']�Z��G@O/;�[3㴙�E��^�g�K\�W�>���MEk�2e����2u�t��p��D^Y�?-%A<iй/���8V)_�l���/���`�-]�����MG����k�L�xDŶ�Rh�۫E����I�e6R?gb�*P�I_�
��F�*��烻g�(���>�½DBy�C�gZ�~�����ef�y��br����d����zҩ|Q���ׂ7}F�B�������Q֌;0b��w�Ws&�t@���11�B�󋝣�Ж97.�����aæJ ~�&��7������>˳��\(�a��T� ��������@{��ϡe�E�Í��M>y!vhcٗN��dN$$�D�lr�. ����Y=5H�Z��[b��]۾3O���7�������4��DЍ�E.�'�V�du!�]�����z�M["ߞ�HfD�cD�pH�(ayP�̔p�����"��%��>)�sbZSHB�m�6��T�qB�o�D��ǲwD-�F(^��F�v�<f&�#��ם�����.2I�bST�؇ә��"M��>:�1�������O�pe`�	�~F�]�W���[ �����Wq	Z�4v'�BuFV�"a�!qz��QN(�iEx-�Kc?�7�X�ׅ�e��m#�4��tĚ�X0wȌ��^ �:Hj�VH�"�(eF��ڐye&�{cX
:�\���<�*�c(�"�U��ւ����˪�+_�G!��  q��rgH�e�PsX�9���kՒ����FzQ~�{8ޔ�^Y.��>��gO�˼�m��� )<�M9Lv��{Eѫ����r0��kNܘ��Q���]hﴣ�U�:G��>��U�&a�gXH�S���;�}X��F���g��9��ఴ���un��"'�i��h��<_Z������{�@�r��a����7��ryq��κN�z��������e���Գ��!M��w�m�S�e�����r�z(�Z�ギ�b�8'/DM{�"o�[*[v��1�J�Z}����
�)�MMt�*�WvV{�q���:tMn��C>i%�xt��;:�`�vN0h��ަ8LZ��<�zƻ�ps���Z����������g�FfN�P�mz�����޷a�g-N:��EqP3���vvPH�]�F�5aN;]��Nyf��rh=�"w{��>�秅���a�Rb����-I3�Ro/� ��\��\���Tl�%/���̻�C��Ab��lB��Bw߰9�����}6.Y�� u�>q�;Yr�h`x�G�|�t�iO���wx4o9̴�b�I #�Z�@�*B]w����}XUd�yӪ	�G ��a�+�we�R��k�$�\�g��'"�t��׍Ҍ�Ƽ��!ԁGx�A"��	�Lw>"W#��7�b[��G��>S��)�(3����)az/4%�Q�T����(��/㔲ښ�!{��6X3�x���v[�]���/|�F�❕\ԃ��<���=�K��s�����
���V�t�.�u"�S:���xw\��"DYrB�>psi1��4�W�{�*����X�3���`��p�������c~�so��N{��cծ�aL������R��{A0]��������kk�~�����n���C��߭4���ь��d�>o:}���`�]b}5�^�:Q3ăM��e�0�@�ϸ�P�C/赋�:!�_�t4���(=H��,�a8̰(�=����s�3��Y�^^�G\�Q+f�n��;Ӡ^�K^��i�6��L�����運�?O��ۊ��u�h�	S�E�w%� ٙyD{՘���X���_���)�"	�d�5&2߉�����0;Յ��O�� �>Ғ���x�#!ֹ��`�އ+��)X�t�ﱼ��.�p8���L������1Fn��җ:>p
8��RW :���wC<��i��(4-n0��~\�a*�u�����a5�Pb��ڮf*BY��5ig\fhC+��c��0�4��C�$����q!cvp״K�`NxW��5Z��+,��2�/.Ī���=I���.�A����>��T�;#�s���~�����Eu��5^�L�Q��Z�0�c �?]�#��GE��$Ċ�$�r�ِ^j�Oz���j:�v�Za����cLV} 4�k=�|�I�����w3Iɉ��[����=�:JMxZmM�M�@�'�N���_�|O(����*|) Q�?�9?mr���5("o~�W��b8���ϩ��Ͼ�8�Iii���-r;QV2�:����L�,��O�Gs�h�zas��M�)S!��MZ�=��'9��b�}!L�s��P߾r���Rǳ��N���0z85,f~�"0z���ݲ�ֱ�o�2^{�qk,8ɍk�}�Ra��y���Ћh� �\C��@�~�KK�[��Qx����/.X�}��X Մ��aF�����R�sqh*ǡ�PB��R�C~�-�$�e7=;a�Y�w��H7	�o�/��DhE�l��J�|ђ?�NM�/qr��5�1����]f�����!#A[�wl��╟�����F7-�W�u�0 _r���y}7 M�o��z!F���ܰ�Ym��1�8�ڤ��Q=�	/�t�E�v�����W���p/�&5X�G�[tI�NΖ��i�y\r���_����W/�!��L{/?\�ȩ�e0�,-�ۭ5�*GL�����=v�=V��j~p6��i�V��µ#sߜ��3��3�
$^�|9�n`�f�X�NY�������GW��|�z��Vd�-Ig��gvݢt�O��ѣN�Q�iHC��q����,��q�z��9��d5-�����ϻ*���M��p��a����<]���#��4.��!;���%�%H���0+���7��k�d�Z\S.�UP���|/xl�`�����ߣw�HL���Xf�+V"��Q��cm�4���V��na��#tj�5 g{��t�C�ߥ������#Ǧ���#��U���4ak!�Z�Dr�O��\�q��x�AT1�}��geL�����g�?#�q/0�20���"�w�49>�/�g�T��:M��p�e������WG��(N�S<�h����iϿw����eyC(���-T�{��\�����r�F`���}�?��6=J�?+�ԲagX�qq*s�z��IM��Ԭx[Nh<@����� ��5��}N-���Ŀ@<�$;"�����Y>���ꮗ|/�̿��p]Uա�g�ȣ��H����Z ��9#�k[�,~	߲^� t�����T�-����M�׍�����v����N�Q �� �q�[�	ge7*Z$L���\��w���:�촦8`tL/��B�}k�[>���YR��T�FŹ�G�#����v�N�!�A�Z����6s1sLS��7���������n����_�ⶉ�wԪ�|�z#�u��=T%�У_1��+u��ŧ+�*�	��3��2?%".(!kk���M�k|g3i�9�4��8�~��?����y9O�m v��`��ֺ��(�2#p=����|�)��)��+�B�j���e�[Xd��vǮ�oZ� L��$�R�x�{���K��t-'�A[/7�!~t�īZM���iD��Uu�$#��ӆ��,�يi�Z�ĪP�v�zW_N/o t'e�a�=�q��d�s����4/�&T�!�ڏY����N+����'��>��|��bqEg'&"�1�J��?�os'��<������=���l�	e[.>��;�NI|'*C��tF��8��(:k�A�kx�<����箷� �#��lJ�K��b�
��Y�[�xY�á����5޾�#�a<�*@{��f�~�@)�����v�攱���=ܯ���&Tʍ�2 �����v�Y�v��֋�Ƀ�#�
�qկ���oa�+O�F��f���T�4"����Ue?�9� 0�U�5��4�EW�'
J���j���{�����?GR�������~��i�Pd����9�FN�C0�֝j
�Z�5z�-�d˄���[�n8j����6��+�.?!��F�1ө��s��*�ӑ:����6
TP���#�pt=�l��v$�S^&�����|�J%э��R.�-`wT#�ha�#`���ݬ���#9��\Q�1��u�x_�m`#�;�*2F��@77d���XZ��p#v'��4o�Qâx*�z]��H����iR�����	�Z�ѿ?
��{`cMؼ8o\�a[o���:�¸>��K�Z	���zqN1u��;%��
=����/����H���bY Ģ2�}��j���y�a��X�#��n��i��ËF��]@O4�)�r���C���D@�c{m�A�r�>n�z �9�h���ƭӑ�UH.%�k�)J��j��U������Io�i�6���#cC�/ٜ(�;j�+]��r=*ݴR��!�;�gc�lQG�`
��o��jKs� ���$��ꋭ��}|��rLk�;.������M��
h��Xq8e$�z�A�rs��.���T��X�1w�9�HXo�D�J�s�0JM��whK��t^��Ș��Ѷ�t��W���R���W��d���-y�%o��?;�䍾Qζ�V�R[��d��`)X�rE<�����rt� �Wl���$��!S2o��7����<�;�v��̓�h��¹���ϐ/��<?%k�}{[��沓���PƮ��?���~�ٳ��m+�$�a�hXڬ%��n����<]-~��D���I4��bD���.��
MdH�6�%)���	�k�Vh��Q��M�bU�y֗�}���3�(�mo4��i���D��~kVU�e�����غ]�`�~��6���qn��?݂l��b
p��ܯ�i
�>��\��:����y�Z�Rz�J%��Q"Uz��XP��k��{��Id����Rf�ઢH��^Q�j.��<C3#������R���֩81������=O��5ҍ�m����u��}/O:I6R +�H�aۙ��*�@�H�h�����M5U�L�Cr�M��T�V�Z�ٯ��\���s�gAx��, �[|�Ҕ�֊@8�a�����t$�kیֲ��Fa�h{> ���֍�4�IͲ�m�]�7[nI��)��8�Ľ��093��U<�����_3/ ��J�i�A5\;���ͽ�\.�w��c�h�¼?�=��-{��iO)�\ս��|q�"L��-c�8�Y������ݛ�J*����hG6��F��z8ҩ6��~CP��k
���k�\忡S
�{������R3�9����#�/Ҽą�+}x)J%�č8kwt���M�7>����P�������ꋟ�WOb�ǙQ��"r�)lB�c��t��ǖ�S��m硙��m��f�	��C�Vl��GC�K���h���pQ�`���6uT��;?��n4�������W��O�fZ�����m�O���
k��/�a���\���.���!��1q�J��%C�����S�O�&������C�Yщ��7p��+E��z��A��E���i�l����)/g\�38�����r�I�,ĝ��:n>fbb��cE��#�=����_��t�n\�Uh�R۔��pt��^)���&9�=�k������D~��ش�xUH�ݣ�F�Z��,I�Cڶ[�Y�Go�4���R��� ���+Lu;}�I
-s�� ��B3�3tg�=m��x�\�p�����,�͎oh�cV}H�lƥ��r�eI�%�J0�r�JjI��A���;箑����|�Zݜ�g[H*V���إ_5`3<�^��MuG��
Eq}�����6([�P�#�Θ��I�5#�ɚyP7P�3 ��@��\
�vci�t�F���C(ï�ކ�G�~��D`�t���� o6{��_�����\l�60�W�t�?�I�K�A�1��s�x���O;"6̽��%���ˤ�dy���QQM�:��n�]Rs�A��R�n!�98[�y�~S&eUv�Lr��~C�n«F�)'��8�o̻�����Z���Y��}��գ���Lc��S���qhv��Dcn~�������D�\��}�X�@c�r��^�m�{��?�V��噅���!���\�O���|��N����j�=���9d���<���+�̴T]���|�8�;fh�j1�]��DOa�J�|��I�>�1lb�O,H�:$\�D������m b�iy�GK~h�ظ)���rbE)j^���Aw� o�E-\�ۙ׃���2)Y軸��1}&��eʥ��５�*dq�>r��+�ly-�'�%t����Wny޻G#��qF�/�
�3ͱP�M�F��w�9U��'J^��}��r����v;Qi'�Q�����z���L׊����9b7t�*1z'8d����D)�i�Aq�|#[��Q�x���P�v�ݸ5Τ���_�\�'�ʱ��u/��o�%5���� �����;`�u�m���m^�Z�)t���H0�S�Y:�`�yWrg~-��+�J���+�|����y}����яb�:9j_��hn�d��+"Ci$�PkqC��agv�Z�@��0����̛��#���'�:y	39���$�U'���ɍB
3j��+�q�I˪*䌏@6f�a?溦�O��{w�z_)��1=u4�O�\����ǵ�N��u�ϻJ�&2(�Y��Se0O�+ʋ�V��,��
������ݡ4������c>��M�Ad�����*rヱ���c1æ<$,�Τ��z2�1�DUz��7��N��,�-��I��!ZBμ�i�����&�S�/]1$��s�ا�l����Ы��3�>�M5�J&-�%�����2?��t�ǘBjQ妟gf�;W��Át����V� ��௼nV�qi^p��^�P���<E�vW:��L]�}G8���W�*�����J!�y�����%u=;���ϑ����7,��VG�B���R/�ד�Q��RUR���[��#���	���8O��!��1C�<vwt��v�����1U�m�$l�jX��-�%Q6=<VP(�<��7�*o�̪���On˅s��7˟T�0��2���p�x�ߐZ�d%~��"liiY�9Z���P�C�@NvmN\�Ir	�n�� ��͍��fӫ�R�j�V�%R+=(��N�i��Q].q�Щ�K5�	�����Z��tG�����)��˶t�4�\O6�	l7Bk�h)���*���.*�I
N2�k7!��Ge�Z��ԡ=܃r*���-[�5��b]~,�E�s&D�}e�a���N�[6��;�4	>\����k���=6�2/b�n�Z�r��f���ITP�u�d8�6oXD�,i�j?2����0�l�SM�D��$~�=b7l�A�������*�Q��J}86����8XD���/�~;��e=x�^�Uwp�fք�!{Ϛ��x�Yl��b����X��	K"�j�E=��~��	ω�3y��_?]쭟^h�G��QC��IC�aFu�u��Id���׷އ�����ab���p��moM���Qw7=�"�^�D�3��`r����g3�-c����Ȟ��\i+�7Cp�D)ݘR:�~��b��N�1�����'�H�2~������,1p���w#��!>M�Ʌ@�o7L'C�$P>4П��>z78���F��>�5�0�	*�퐷�p�&g>#q��F>�SQí�^���\��|��|����lsT��]'�����v��W?m�����E��v܍:�������}}
��݇��Xg?�Z��?�<��UP=�#�x1j�JE�W����!�(�Z��ax$I1\����dU�q)�麕��0�2�=^��aB$}������<d�Y�������o
v�t0�l����E��c�U�.0�M��~^�^	�W�5V�{vc���_���0a�M��xq:�F�)�_"3J.�/|i�y�y����~E�;X��K�$�
��daL�cƫ&�ʷ|O(����Ʉ�P&���l����l���w	�
Q�5h7y���S6�'�%�Y]�O[/����Om:?W\�5AV�{�i����"�~C��Eq,�<3^iJ�v�M�����\%���L�"�n�5�{jnaf'���L�=u$N+K0t ��*|h�2f�G?�9�$�ӅWS c�����R�&| 6�]���c&��	�U��G��p5i��.	5e�9*���PVkf��p3۾2:�	3��,J���c��Ț��n*���嘒��͐�1��aކz�]%H��q�37�:@�v�<�m�9������*W�'�=�{�gs�IZ,���>9�^@�߯��^�+�Γp�0CXn�I������B�[�#�q���O�����ץ0��ٮ=�y��<_d��uݯ���t����>�^_<P�e?^����#�P��K3Q��2`z�A��7�8an��`-o�j�a�N���~wB|�7�P��Z	8�!���/���{�;��շ�B-�V�׻y��x�<5��������*D���C����Wt��P�`񻴡07=�pn���H��ܝ���ÔC�w�1:����Aڼ��-F���o�7u`��I�^�_�j����ݪ�&��B~T�=���C���*P`��av ��J��a[���VJ�e��V���a1�{  �B��w�U���Lo�����Y,��f�X��NJ�#猞&��}Ч�&#�k�C�Ͼ��g6�G��ބ�S;R΀=����e���[D�ǹ{*��"rؐ~�n�8B�T_�-b����:��3[��Q*�|�E��li�(��}.���U��o�@/�m��*&����&&�-N�.;�Y�w;>��
��vL��@K=9���	1�סchV���-�6������we�,&��~���K��<:F"3���Q��]u��	<��C>��h�����f ����x(��[4[�5�$���՟&6�G�&����;���ª�/�TQ;9�X>R�B����!)r��^��ђ�����7C���]z��R��i���i�\�
�{�B.�N�_:r�ˣGӄ��
���xR���cF�'T�CQm-ck��GyY�xN��+�.)S�oCƦ��u��Β�hEgmǫP��L�s�����]�,3�d�`=x�����5,d� ��7�i߄�f��νϵ��An4�2_��s�T�R+x|_Bp�D�g�B���!6�G΢ou�'�R���w�B����ԙ��z���:7�Q�5�]�K�Y�w����'�l_��bj�O��"�t�vj�_�L��ڟz���+�M��cK��.z��A}.��ߔ�� o�6����J�娽�&Ȝ����D8]�+◤����O�KS챔�^%|�U
ִ�PDs�vw�)�����ל˿��
��ZM��E��:�2�`/g|�#�WRS3"盚5�%�<n'T���欑:�y˩F%�\�%w��M�wԃ:�j��Tmt��������67Y�&��G8��X�!OW�1�E�W�r,�Ge�C}8�l�Xb)����z�D)�$ lqښ��a�M�%�#}��h6c�,̀yD� �⋫f�W:�*��ڂ�}���ŀ���K��C?���GT,*2f��!���7f�o��B_���FWҥ��?G&����}O�G�����zqL���&��P�O�����7��C%Yr캒o�o�����:ϔn��64q�K:]�E }���9_]�Q0{D��@�w��NCq.\��TGNŬ	��Җ-�~]�5H3mq�O�@��t:Kl�f7����A�A����~�g|X�oxk+]!�����I�Ir%D� 8�8�V)i�ri΍������<H-ĸw�h(���U�$��?B��ÏY4/��������]��d�ϑj��94�n����i�*Y�~*�����«S�ė�&ASx�e�Ã�'XY��.-��n��+&�+�ى6����}Q���|>=�I�W����7���w'��IR�JsΘ�T!�2z�(��"���7zDXT{U�Či^!jyy����`_�_�L�ib#M��2Ԇ��&sYE'���9��d���c�Kk��Q�*8���{���,M�u��W�)U��i6U�S�����_��5�:��삄7�f� _�[\
}㞟�On�O�O
^+���tl�����!��n�]����!�uP�ܶ��?�<��{o@I�ò����^��d�q��dŬm��=n^P���d���;��G��8�p���h���-K��� ��Թ����L��T(��G��F��b�!�22>1,�wCƉ�����v�N��ܝ-#�"�߶�c��/��h�en�8�J+=���D=�?]�H�n8oԥp�	�����y��CN�_���8zZ�9��p��"����L�j_��uĿA 	%t��B1��7aZZ�S|����c����oj���&��Wſ�gAA(+!fp�łT���F��5Ǘ#��O����������?p���	��
2��������_�=�E���M�C�{}�Q���4��/PK   �8Zj˳���  )�  /   images/c68186f3-7e1e-40af-a8fa-ebb36c358ae9.png$[T����0a�2���� R�#FH�#�;��K@�0R��n�����ζs�{����g_4�p_�  %EYm  �3򙈍��D�����M[AP9F��|�n#�& ���=�a ��8+~p ��=Q�J,��N%Y)]��^�/go��3l�9��ڂ�y�L�W��g����_��0�|3ȯ��?�80������q��2�����srb-޹O�}�����B�[���ߊt,��.�;������[�w�:��8��g����ftk�wk������u�-�k�	}:���ek���3�������{+����W�=�2����4)%eT�pj��0%rG���D��G��Fk�q|l?������# ���R*)�k<z�븄p��d�B:��  *�E�z!����M@�u��`tqEq���UT�D�7`ُ�XW����#�p�A/�VRS��FH�`�vr2}+��fM��DO�ǇT����  h��;~n��$�"ά���Z5򙑾����(H���ǂ�����������Ii�б��^����Ž?lo^�DN���?2d�C^���*D����7���}~�y\�;����<9���z)�)�M��.w̅�R��Q$Ǆ��AxZ0�U���X���� I.�k�~k�S�,��7lzIT�,m�^�C1�XPXXx[c1�t�J��gl���`������d���rs׻���>�h<\��	���"�a��Ią9����#�
�O��T��z���\�`�t��.:tV��tvЍ�A��;�61jn�XHv U��^kHHV!�,j�F7�����F��q�`L@�F�8�'|·o�mG�u�_�I����ֻ���0.y��.RQ$ѷ�8����dz�O%��-@	T1w�)#�8�eff��==|�|�!`�2���t�@��t��������X�r|�*�V~S�qsK#��R��n'����IF
���&� 3�?u����(����s�b���NG_�X-\�B +}D�P�;��c�נ� M�6���o89*O�ᾫm(�pR}�N���|ҭ�׊)zxhh��"��L���&�7�d����c��-�������q[��Tuќ=^�^�o��j�����5���IЖ������ems�s@�dz�{��u�Vid�ģq�c�<�Ȟ����*#�t�a��6.�\eP������Gw��X��R�	8����}C�ӆ,�
���F���6��9�[�oJ�gI+ӉckR؍��8�GW��+�g���,8֥A<����B�
wd�ۨ#�4Lޏ>����K�7n�ؖ���,���]#|�I�A�:��g�6��>%�	�o��6G�**+s�!��pz��h2^�,����F�7��կ�s���,��W���B��.g_a�|���"#q�vo-�N+!S��:�G��ǶC�;"@z�}���0�n�Q�q���,߽R����2�W��j$�E(�����>��d���b��S�'|����Y��t���74D��K<t+��\��G�������ee9�^cM�Ao99�+����k���Ê ��/	� ����*���������Oj�k��qy�/)��̛EĊ�|�:�W=�@s�[W�:JKo�V��ɮW�V	�œss��8j�	��R,a/
x}�"��;w�;ڋZ�
�_�3!�7;jd;x�&��%���!cLHW���3�����c���z���n���L=��YE{�q
�R��t�j�00R�5��.L0\|�a�JV����F���)Ũ�u�������^��j��O��\���1kQDy���yPKG�����Į�-��>z;]-�,��2��u��A��#h	�`ҽ�Ϟ�dee��j�,�ʅ��EӴ��3%��c�r7����-X:���]/�]#s	YY�0fHT�����e�=;s�r�EO��6&䕜��A�Oh����ʶ���.��Om'�1�I����hR�"���_d�&��<">E�5΃�[#inc/�.�������6@��:� #x�#B�/LG\	aN�,�i��'LI�����U�{��ʈ!��ׯȍ��載�w�
��U�UF)�����Ǘ�]����V��rs��+2�As�s�6�&}'|N���<�2�l�n]s�#�,=�ն�a�e(�?g\�W࿼�(�g#ۛ��gg]���^�s��G��Δ���y(r�X^�R���p<���)ZU��/���լ���@�8�Zak{d�p7�����録ת))�N`"V6�egt��W� g�Y�&T�������+�E�dQ�'�o<Uwo	Ky&	�+ :�'31�z$��/,R��/��[D楧���0��8�s(����n.L�/�����B��E���WӔCIEU��4����-�ն[Dy}��r���H,��p�`�?�~��������H�.��(ݺ�v����������`V����*�эԺ��%���A���8��A�Q�'qw=([6B2�D_�f%���w���^g�e!'9ע�TK?#����E�0�y�"��P��K�o,�辽Qk�9��d:"XX�xe"l�s�	S����Ju�W<�+�c���qb�,�r_�,�݉8�tDsx9<]!>*�Gļ�G¤D�Z�a� �6b|`�	�d�,*Y�KR�y�,"ӛ�)-Iqj؊K$�Xrk~�k� �!��>��� �%±�y��F����U,��$^Zݞ�U0�-���-5dM
vl�L�?5-���?����_���L[w����<�lh��Ù�Dֿ+��\<���7�e�v��]?mQ~nLS}h�|�M+�� �4�����n���P���Dm-
�z)��w�!g�������B�[�Cc�pQ���o�����0OߊP�K	�����X�P]��P{���@��7�o|\X��|#���sHD�z�Sup/�,$�jWb9`\l����d��):.3W#5������Ey�9��X]��L2h��'���x�oZ��?\/��e=��K���D��)�O����
�߁�%&�o�۔�<��=~�e��c$�C�Q,����p��J���䣎�)��:��NEl��(�"�5�6��AG?����f��`�FH�*���Cc1�d��F=J5�QB� ���hkrzWBx�[��+�%��),� ��e"���%��ޞ��Il���脜�h)��Y�|�v�K�I�2.��WD�3���5#�%��'�1{�+�l�])���zAE��[40(!��r�a�����:���q�j���rJ9]�/�z$:��Z�8`a��u�5�ː�tw��Y0jѡ7��i{�)��;�4�<)`8�����4��ނn���"��R��+1( M{�y���±zyBj��>����Ҹ8��ג~���:�7�Q*TRyv���(L;7��!���:��PN�_׋0�Υ�T�Z&Y��GO�!uU��Pq��޾#�0��$_�'}Kw� ���������q��?9_d�U���3G�t����	�eu�3c�����_��`W�0��J;]&��f1l�*��ēG3��H�ƀ��,aeUeI����\��l:�j�3��cZS[g/��.���?�!��</�������T��W�3t@�e�%A8�]�h�?�d��p��.o�y��L,e�g؅��ټ����O����k��À���R)|;jݯD���΅�0)��󢒄��D#M��ˍ���	cq�玦�E��K�ס�^��*[�H���-�~�����n�[����L UD���T���E�����<C�S��i�Χ�M���xly�Ҷ��\�^�hx�2Y�䥌l�(��6p:�����a�Qױ��Ε�s�jp�ݬ��G�����0�ױ�=!ee'�Dee�?#_��z�?RX��Q:���ޕ�L����lߡ ���������`�9zx�h<�����Gx�]�������?#�A�v2���8�YA�_?�7sN�xG�[�5-C��6�l�~�Ӝ��G�81b�n]��^������M���$'\����	�L%�� �~a����jG*�P˳�;�"C����Bw%�Y��CX�͍���2)�z�����q�o}��5$/��<No��~�2�U�Y�G����� �5Zͅ�F>y\;n���;��-\�(��@��f��ՙ��{l\�?��G-�"�m	�s�3��c6Y� W�Yp��rq�%y����T�^���9�v�1j�{�����'rTy(553�>�5H{o��d�)�.H��fF��ֶ�W"C���N~� ?o��� �̔�p C�vb�r���r�p�AX��;P��7�R����-ǝ7�&Ɨm�:<��D�ت�0*�%ڀ��t�ml��
�u(�X3oN^I��M�w�f�I�쫪9�*�d��DM)3��T��L�ѕ�J�8C�cDmEf�����X*w�rO��`\�ׯě�>14b�s�D�7u���s��6�)���֡$4 i0�Nz��"��8�wQ!���:`1Q�r��t!����j�% ��b���>��R	��'�n�M�����j�y?�ކ�EG��KuQ����u{)�8�Hn%��ξ�)����1Y�;�Rߓ��S��������J����񃅺r����ߦ�܅ ��x©+��!U�o*�:r���H��Y�`&ƙ�U�(I��CY���S*D���l��h=s�����E�9�9;��B�OL�P+
�	�$�����p㐲��Fɞ���̪�'���b�����n��g�3N|Q�JQ���v��q��8z�>[u����γ��܏�j>�7߂�}�������	=H@7e�`�e�S��}�~�˪��1n��>�d�Γ��Y�w��l�ڰ1������s�A�+�Ȑ�5Վ�$.
�^H�����
b7�o�)�+�%~d��Cn���4Xm��0>�c1������Q���b{t���K��)�̀2k�@l+�B��vo�B�����V=��@ig�m��Rb�<c�5�Cb受���%��������m\c��7{����M��V�m�XRR�>wn~�w�N�w���
gBa�e�(%^�1�[��^B[��h�?��������̍��`3���&�TD<��TI�.�i(z0�l/s�ʾ��03Nh+5>��a�䄝@�0}�32�q�����]q���v�9�XE�6#�ǣ��������� Y;ɏ�w�l�[󸬗��������{G`�8�q�sv�j�'À��I-�wMY�E��GY5jo#9���nh�h͌����'{����uEL�|-��f���\;ԓ�py���n�5��<��p#���}�"�8@��ޥ�{[��
�q�{�w��?�_!������t�����}�*����������U��B7�AF(V/Ƞ2(������x�|>��X6��F�>��H<���X�����sTe�X��$�.�����6rxc�����wr�j��g�N���CCʮN��[+����� �H{��G��H�u�7��ಝ'����j�i���\c�jv����Y~���Ǵ��B���#AM��>
6�/[��"kO~�j����T�x����Ϋ���g�fb�H��"`�RX��/
������B���l6c>�8��V���n1"me�H���b�'A�#����{Ī|v���!���K����CA�BPT���q���ެ�.��h� ���{����T��d�D.Oq*�H�9�?�>9���s���A�g�S���&̪�j��o�"��zo�$i��tE[�*���o�Uz����yD
\���۷]T�Φ�X�ndzZ���Κ򜐧v��P����*����N�$�]2rm��Α�jW�����dԨ!�Z�O��HV�0f}�R���3�-������� ��S�#����4.�|2��
qР�~��vC;mk�&5%Ts! h"u4�$[Њ�!��#�ü0�c�xǳ��X�	�R�GN�$-�'ZC��.�P�������xd��0駬R���9�j��Kп���f�]����l���Åy{ɴ�%7�������dRFbO��ܗ�VI�O>�bW7$(ޓ���i���#>�5�v�|a�!8���<պV�>�VUWB�P�9��B�M����ft�xs�WFZ Gu��)��ʚ������SU�;�����O�o������%yA��lý�M˞��Q��Kxc}h
Ii>00:�a���>b/�䦶j/�NzH{���s|�q���ٗ���\S	��`���r��W���g�;��!@��A	qge�F]��i  �NGW�4z��/;�\�)Hd�b��~gq�|.�¤���:i&�2H�w���p���oo~T^�)����ʲi���C�J%�k�b5�O�Ѱ��"���z�Oa��:��c�[)4�ubyFK{�V�/M����>�I��s��i��U��_6OD!�c��$TǏ�����ӊIGs~v�F̓��Y����ߦ�R~l7����ohhPY�MD�91�4��|�"x?"Ҧ=�v�"�r��5��Ր���?�G�;���~c�<��;*�qHw���E�������7�@��@OI��@�r���7��e'�(k�**�G�%x(�~L��X�+��`��� �U� �!z
��0�2�C��m�r֒�S���NƲ"�CIU�nW�|4X#�F�붬鑒:ܡ}���l��i?�����&�
Uֈ_b P.E-�R8^�S5���u���w��-�h~�Z�0��+:j���Of� 
����E�,_���)Z���Pp�iL�!���`���?Ī__��'�Z�� 5�x��඘��W�^����ŷx�^��	�X&|U�!/k�B�9'��%m�zc�>�RX��ƽmV
�r��QL�$���+�]4�:y?���񿬨c-��\F���o��b[%^XS�e܆�LIf��{Ơ��n����i�c�Ρ��:N��|�O��q�5�_�«ܘLF�t��w���"���k�m@�.�V�I51h�4��G���@mLŏo�^NN.;^���ov�N�E$�Cf�us��qc�3�}�+�檹ɕ���T���W�u,�e75Y�-���x�WV#al~{�E>�68���66ě?��L	�k�OJLnͧg�_�������|)�Ab85�r���
��M���_j,?������Qf�罃J�ۗ���	�$�?�ԙ}	�{[��r�����w��F!h��4*OR��r��D���:�gp��%v�ϓK�n�8C0�e�3�K��|��qrN�������'�u�h��D�X&�㞓����g�����D2��y>���D�G�.==fEh|�?l���L6hn�C��~�q�e݀_��޶����D�e�q ٲ��f���l������x��;��L��$�/�eY]�t��t�g� �"����%�LY�j�Z0��\�.��}��9�6.�s�pY�ە���(S�l�~LK���!�0 u\���g�B$������=�w��ڑ��,J����������а��w��t�50�"1���ȡW��I':|�{�8D�,��n��1�dRqO���WA\G�8���v��7J�n�R�݅	]L���2�o�:<Ufĭ�^�]���n��7	���oU,ԖL�w^(Lyz���$�:j�)޶5�?��bk���� �H�x��_
�3},Y̠��;�>+��JN#��#M0��)��#�޵q���*I!�P��Y�q�@�����7h,L���N����s?٦/�?{;^���W�.MLh�} �Q������x��J�R/z�4�n?�,�}ix�P�]�6��'��{d�םr!�w=��Y��-��t>:���曣x"���P�n���%����T�9�� �"����1����A�?C�+��k�[�+ٮc/ø����E����f��'�+�V��Ţ���]�N2",S��9��:r���Sނ6�x����W�
ω�0HP�	ͪӢ��^w����?7���>��	m1���?�>Ŗv�3*`"ҩ☒���� h��v�鞶�;�<eУ�<xCPp���R��YF�~6���l���0����E,+���2��!��H�Q|���(�����1Q�V'��nu\�����&���Q!;�.�|���� ���@zT9��%�1��\X�ȞQ�-����r}��H��[f6U��Ԙ㆑�v}W8�LA�r���r�<����릎�������z/�Z@��1]�G���,��m~ӸM�/ղL�zgaѣ���P��f\����|#2�o?x����4*��\Tp)tX�����S�ti�;�-<Ox�ByQX�%�,+��Å�;��Ys3?t6�R��;�3�	�=�+(�ͨ���%�4+Hܡ��ut���vSX~*��T������_�vu�|�΄L��>���s`=`����k���Np�'IU�b��_=x��ƬҢK7)��9��֗�G����?���]�O[,�$��$i������~k39��ϧ��qu�p�w�3YT���,U�oM岐��NeR7������x��l�7
ӭq���+��}�#����~2�W��V$q�5:6�p2q����^J���U3�d]{#���ĳ���+���5��GD;;��64W�ݿ�!ɰ�jўƙ�X���������)}~��ߠN�ϻ� Y�%�6}-�!M��\� �4� �O%u�HT�r7Wo�ko/��4X.������ة�����[��1I���cC5�@�˺N�3*&���i�l0�v�gF�ɣ�ܑ6��W����W��G��>R��o}wj)�#�ES����s���v���ۻ�Yn��3.���Nǽ'q�1Q���x�ݶ��%x-b]׿�ߺ�n��.XFX�,%�=Psp��۠��8��r�j_����Z(ai����{q�s�ȵGGG� ����>q�\�gw�|�`D�`�T$��MB�ߡ��� ���A>����.AH�����mo{��"Vg�c�R��'�Z�1Ly�kZ�UA��|,������vU=�+|w��:C�4��]�������F-�J�
v�{[���10���,�y��K=�4�V�8 �$��1�BD�1#^t>u��_U�v�����H	�F[��p��r�7�i.�*���;�Z]�ׅP����g��>��ȵ9��b}��+(���ˀ�^����"���m&0���殟���܍��,�RjY��|5�@���$�W&�@��u�a� 5?֙��dh�ו5�x��DQ�8�_-�~m�'�Й��g���
����}F����������6U�~�v�۸ص�ڴ�W%i��-�"<K|j�A��Ü�7�g)d�С�&��*G����d�ˣ�&��6R$����<j����c�8�-�eU����,~5o�/wh1�����G]�O5���R,�f�1��}����23b��
�W?�)
���҃^+Вi�-��x�^�Eו�^	a����0��n��i�L �z\��b��a�̹e���`��v���ar��bȠ����L2�Ƿ�X�\�aH쿘�����(/yd��}<*�j{CPRI0�O��2���b��#R��;R���ݞ�ƅJ��T�$�(�|H�����cjl�=���*������ ��#�+W�im�j�,2�{���	^h�9��v�,�FK�S����i<u�R	,�ϦW�i�$�2:}����o3S(�5}b"�)A�@K�1r듽�Թ�ټqC���������a��d������_�k���lƳ�->�: �?x.�l,��	�]�=�PҨ�Ӎ������9&~���Q�e.,��'4���$��@�v���11��"�ۑ[ l獖��M�����i:.;�^c�2��c3�!���ls:H�^X�<UZ�b͗L九Yx
%A���n,u�8���R�<aٶ#rU�*{h�h�K�y�K���� RU�I��N��5���$������A&��p4��D��ʶgg���E�.x4�b�K��,���h^{{Ѫ'�0�0�r���d�� �E_���K&���hͤy�J�D�P[d�C��*!Ik� C��xQ�洺2>77����h�w�a�]���)ÇH��E�b(�@õ�����譕#<���Q%�D`�g���«�Ү8���Iy������bv4uy�"k�k��g]e!�F��5
��,�����>��Q΄�T�y�V���L�!;�:O$}՚B��e������ͺk�>������L;��_��g�VY��=T�uͣ���o�o��Z��G>��%��8!��8�ې�i�<���S�i&/1Ne�(�oB���8�#�!p�+3bkk�z,�Æ ���98�ƨ
?j�<aa�_�Yo�d#b��a��dځ̛���+R��N�����Y4��
X�4M �fģ��:�KN]ztb�@Tv#^�6�֋����t�#����*����;#1�tB6��
֒�jOd��Q���qX��gМ�����h��&�1d��C�v�����&jGo��D��ҫ����SsK�0�YR�B���FJ���p�E�GAƋF�m��F��W����������
��z��گ��ͷ��:ؐ���<�f8�Զ|�Z*K��m3��-~L�j�P��>�m��!C��r#t9A�� ݡA6����G�x�o�������u�\��\�׳5��d!�◫����(�nk.XF��H�~8ŗ�@��HL��v���7w�3%�m��m5��M[j�7s�)E���J
i�G����������>y���h��+��]��5��?�g~$D��X���V���h�=�#��9������QMS�L��/Pv#��5��s_������rvQ�84�� Ӓ�>"	���`$ೊ?��e�u2�=yZY~�W ��6h�Z% ��߲�̄��0�'&�JTy6OK|Fޫ�����Oꈩ���g�)�W���ǧ+��9 ŕ~��e���M���P�w\ �vv�9A5�6�Ẽ��E=ƐJ��Ϗ�v��uӨ������R������7����#a�g���p�n��`�)��������3f�D��73�ׁ�6�sk�&��-l5���*Cz�.���WW�������慆��>���dĘ�!GJD%�&7/g�
��������z&u��<�e��v@i:zQ���3�.C{xW(���иGO	��V����F��A/�/am�:�C�U�� (Pp	-B^i\������ZY"�{}�$�{m�	<O�_���&��)�r���	�RV9@IV4�k���A�8>���yU��`�U�$K����!(�N��G�c_U�<��_Jqa"C�~gw�伳��B6K��C��wX��S8 PH���8��Ǹa.L����J�yY��cˮ�"��[꼫�J�4�Y@I�e-0�~�Ά��/���U�nB4�A��܉ӎY��j�Ch'>n+���+7�Ca�������F<���!с��%?>襰�ӡk�R���	�(�;n�o��*��4AU�w{\Z�TZb<�my�ւјaѪ�Ϛ��H��`��^=3P�?o�)t?h�,D�8�Vd8#��H�q��<���Z煮̫��*��N@�@�+�r֕R���������v�hC��$��򪫺��w�M7䆲&� q4��\~�gK��w��j ��UFP~b�?p��.��%	I�{�v���/[�"SnvI!��&���&3�!n#\Y��}�"��Kt�O�����č̥y�+�'��y$]��?b��M{--����q� �<Nj^����o��Eu���e..�L���ѐ�M��2)g�Vf��e"��E���T/#�w[��Nk��~UA����Y]��qB�*z���3n�V;EC�������/�҉<�cA����q|D��}����:Yۖ��{�r��*�C���p*��R��{up�� ��4�3GB疡�1uC�4�f�����Lĺ��@l��[<�p�B����JM^���EùES;���r����,.�O�)�E}nF�r����QӅ��(�ί��[�u���D����X��:��J*/��-���e���&�o�_Tb)c��a4w��ޫ�\aak	����q���2K�	ʓ)-q��;�*�QIߩ;��1&�
0�u���c��w�8�?�t|����xP����iX�7����~8�r�`@Ԭm��C`Cl�wJ���
N(�5�3<F��pZ�V�tx\�!�uU���ֈq�q�n\n��`h��+�O�ov����id�'1�sa�iѵm���J�$%�}�{��v{L�>�I�7�(�
@|"�w�Ȟ�F9��/��5%A)j���Ǭ!�e��uvvFDзVd+��Z\?]5�]�\�^��Ue��L�S�^���N��s@�������dC��m�<{�!�="Y�C�D&B�_ܗ]l���g�0w�M\xcb���/-�V��S�~+P��W�s`"y��mx�ˎj�ϋ�r,C�s@;x[�_���Όl~ͮ� �aa�$S�`�璙��uGi�Mu��ae�QFo���Y����U��8܃��QFo�|ǩ'$L�����GP����X�YXʶ5��T����%���g�cU��a �0!�0�m�1o^d�������t�e�w��p`*8~{3hy���& 9���=ՆkP��Łd���w\��Ts����𭬬�mߜ���Ƌ��P��������r�'��3n)L�Uq�7l�5�GlxO�C?�q�Wq������-�Ni�n���%~�e\6;��T�;��ؔY�V�G��3�LF��Q8���F��T�Vk��g������$|�_>0?�)���������ѮZ��\��W���-�E�f���cOJ�S"K�m�;U(�&)=�3�|<��`:r�<����''CE_y������7_�m~Oo����vSƠbb��e��}G�:���l�`��gbBˡY��i
f��/@�A��}ggE�=�s4�$�&��²��k;#�P����r��rt
�;�ś������}h�U�4�E��Y��N׶P����r=0�?οY#�ھ��C,T��Ѥ�s�X��Y��bO-dDWlx��  R^��t�*�(��1����]�h�j���N@���|L�al�mk��>Ϋ�zݑFj{��ۿWH�B�B������ D-+�e��e�t�i#�a�~/�W¨���A,���ITL2�ch�.:��r���̋d����H���zV���E;Ł�������m��(p�S��%0Y��D{m�(��^`��ą2��W�::]�<~]Bk��(7���{�߷�7rqI��"b&r�	*�gt1�;L{<�W�G�:�A��(镦r2�n+vm���|����X��j00�r'�ޞ���g��ۗ���ݼ/	_(�g��~>�sw�=�c	����J��c�v�廗Q��'�꒢�>U���//�@UM���?��S`5fG�D_0�U��z���}�l	�u�x��kZ!�ݶ>dtQי)u��S�JT��5�$��NM<������0�Sw|h����?�$��43J�-eF�K<:ңI�b�H��YN�򑭤na�b�\�HEE\����{��TѲ�ŵwP;̾ad��b�-�,��kk@Kk#�����rM�M˦�I�	c?"��GQ�!P��FNP.�r�$�M������B�.WB.9�(P�,�Eq���kM��mR&$q&���j��@���q���F`��f�^����^�1�y�j6{�iޤ��+�/��,v�V��y88Ih?I4y�+����+?)w=U���h��`�R�z]9�J<�i_\�>�����Mk�cv��}D�<'ʝyv��VƧ�4G�\��8"Q��`[
+X�+)��F�JM4,�!���1g�&D1Xv>��uJ�������<���b�'�o�X]��;K̄
�YGv���b�z?9��Ѿ���(`Y&�(/Ý��䳼io��(fo���$ �^
N�b�� �(����Ҵ�´��H	��M4��%`��t�/r�J�ӧo���mD	w�5y%���`���/rk���B�ϼT�1F�(�4�T�	]/��d^�p���<j�������ԍ�b��۵����,\���}�����4�VN;���WGv�o�F� ���<׉E�.�B8�U��)5@������c�:b���>>�c��Fr����Pm��<)G�v�_Z�j@,қ�lE�j����}�����q�鬾I��L������>�q�165{*���L��O�go'f�o.oᩱ�(pjlELyC�$!�P=���9_v��OI5��}ޯ$�t#Ŏ�%ųi��P6����{�w߻Y����EQǠzM?�B�{V�:"Ԓ�6DG=����-��ڡ�h�ހ!bȃlԽ}J̰,��gS���e:M�1�XۏT�
4�D v���	vwT��O�O�98,�-��Yỻ2:�&�엢�֍旓p$;��;�93U0wc���ܼ<�ئ̼wm�6L�sN{|A;H'F���5J4TN8���w���Tg4�d{}�*Kۀ����P��tD�W�@Ώ�X���0���&&���H���QB4˛���N���W�n� =E�/e�J݅+p_[d�џbMᤊZ�>W��ײ���"{�A���߼ޯ�q+��+w�1ϵ�K�\J%ɂa�BR����%��S�j��=a��f�z��1p��QT�9�;+b��}N��AC�&7��E�cڭj������W�M���!}��8���Oα(g�ݽ�"ܠY ݾ���-�:�+Nr����:(� ���A�;-��F�א5�LG����b���d�}!QQQh���M�-��QoLο�ӑ�ۦ˧j_�� �V�K�A�Xh(�݅P]�o�Wej̗�͟�iޏW��9��:�.���1����a���
��\�F��0�|/��4�D�(�W3jI��#�Y��Փ��
�
��U���p(��swWb�JkU|��@HZJ�q����@J�L�1����z�o_B��xՒڲ�|����Л���P�v"6���3�F3����61����=L�eLh{��N_y�e�b+�"4N�n�;-ưZ��|�j���Mz�z(4)���шD��,~ B0�0c�E�&�s%ݍ�ن��o�s�[%�Dv��:5�TB�%e�T����%����v��܏�og�]}Ytb���z��ǎF!H��e>��I-� ��9��1LX&�)��
Kg� E�{��x��I7Z���F���������RbUd4>�O}9�E�U�F���Y���ë"�3ܒ�*�`z��5���~�䪒g���t9��*�:��ڨ������"�~���¥��v�N.6>����U���764�9�S�zŝ�M�^�s.�)�*��(�L�."UPVfWd������z��J,��*�����K$\M�m黐��(��Jy,��޽_Y�ܴ"���a̩L_(q)?n	�~���)r�����	�g���'_+����Ѿz�f�^����_���D�,�}��;����Dśw�x�z݅A-��d�2N�w�Yxe��,k8�(8�;Dq6�4!hҀ,�s n�Kw6g������}c7��Ob�5�N[�Y�V���Y�/��N�Ε��LC��8�ޠ*q�8''3�,����<������8�E_��Y{�%?_k���+�/{#�n�ē�������{�D�}��^��n!,���&p\'�U���J�jG��=*i��w�0���!�h�k>7�k'����؜�(=R�d��pshZn<��Ԋ�*�q��u�%I��~����	[�4�!K8��b�
:���N0�����=�����|��HAК�?�s*h�Y	V>�~O��͔�<�Ο�	���D��F<w>"�}���S�]J���Q�� ����՗��O�j���z/��D�m�a���%�x�/�?J�Jra�����;5�vdr���Ĳ���Y��D�~G�& ��.w�jPKEE�+�(1�Ǻ �e�4+�@)Rz�cH�G�#8J�?�q���?A��?<�^/<�ii����8��_�~j-ĔƆ��0�N��ӓώ��Q|��ٸ�[
#�[v^�� ��y���7wg�ndzi)Y�>NM�С!e����o��Fs�u�]��xz�r�^mZ���U-���sܺ?f��a�$��X� �^^l���R4�Kqp��*�8���-r[T�K�b��P:�qn�t((��[�m�ؼ�[�i��� ��h�:">��a�()-�y�?6q$��6#�Y� �xpVd��rh��3J�،E*.t~���Aq�/k̠՝%��H��i��7����1(�;�?O��kh�ã�i�$ʼr�ihB�����'6õգ���s�5���yT���O2D����ءn�dҌ��is����L���J���W�{���1|����UWNE8�A��88�x��6�/�/�E���"z�Nt!z��uW�A�z-QB�� ZD���������e�<�9�33����k_g��Mf��x��ٔ�j܎3������,��Ǐd�P{�����e�\�����qy���������ZH^��| PeG�����zj��c���g���� �n�Rz��d�t��<SB} �ҽW�ABE#.O�l�����8��7yd�5��I,I�w���=�)�Z�>>�uL�aF��MuX��Sx�G���Yc#�c�t������������g0햀5e����D	����I���V�K�}���C��/ى<�'[�٫�ޢ��2�z�u��ͨy�e{e�'�,��W��tOo{��Q9R(Z�=������4�����j�M�&E�V�̂��J��k��'�-m���S�D�ZS�t���Y��"�A�v�c���lg�n�����i�]�朡�!�����ޜ��7��bd�r=p���r�<��o/"tb�8Q�;Ҙ�D��q��r+�H3_�y%�`ŏ���e����>�p�{[�������.Rxڏv���^�7�+8	�ey3��^���P�1i���m�#!z$�ghww�Q��5�e����T|/.������/ z���n��aTk�AMM-��UbK�\�K�݌���8�*��z��%}@�#��|����UA����3�넦{��D>��&�B�
���N�� Z ��W�a�)����H]|��=6�̣�����ʓEm�;[*�:��Ԉ����!����ka����������K��q���gjqK�L�֣6���`��Z�N̅�ӑ^�Ȋ
Ժ( HZ0��B��Nы�Ւ����zBoY	���.� ����Lxܩ��^�Uq�����Fr$���v�q{!�u+/@:k���/|f����?%O�2yL#��L�� �����T��:�~� �e3�j�,�Hbf�'.-G���廢ǣ���Mv���/��nQ V�d�
�u���~��h(f�c5�=��O�D],�l=ܠ�oN�&X��(��g��i��uTEeeS�_�f�._�ؠ-A����Bu�Gx$��F[�G�i*������.u��~�
�\xjj�ZJQt�?�Zݚ������:�I��?EG��_�(Ѐ�SX��.��j��qGO�m�g�Нɲ"4�)���R�),0U��X��Ub*��A[.c5ґp�~�sI�X2,o���~�$G���� ƺ�Ւ��^E��������6���V߫��mȍ�a��n9`�6�N���=����{���K+*��_(�)X��	�AX`�����ݧ��U>0Y�;�$�-5w�DAǓ� �|��Y��T�ܫ#��k�ߪGK��6��ؙ�aHd��K �����֣�V~�� �ccFT�:�1�w������LF`���"_���bM5y���ʋ�c��Dvx��3Y���^�{�ƸN�B�.	x�m��ĬL����NC�>K��&�w)d��_(�w��!����&Yn.o� �O[}�0:n#�zsp\�<"�[��gѻi_[��O�$�����v����亴��qۻ���:�4�s2_�dx|�>
�L6lPKŧ�yД7ZCA�Va-D�B�%b@�������0����1��?F���x��.'C<�^Y�%'V�P`���a�X�>��W{;�G��E�
ip�{�(J�/�"�-�i���[�f����0��p��vx� 9��o�d( ��oh������z
���J���X/IC��h���f��Y�GA�_��ov��~����ҫ��Ȯ����
מ0R%��A��#f�O����F���t�'t���?v;&D�`,0���S��!\e���9$�O"EYo��l��P������I?ý�/�8=~{�Z_�M���|�Օ]Ct��������1p3^6����}u?�%���qCa:%Yeg�Wb���&}z^���t��i~�nE��I/�:�W&��?7������z	;Y�_�s��=Z����[���K0���7y�&j�T�}(VU}�D���w6}7"W������4�Ʒ8��6��P��\}5+��찱q�;����i0)d+��q�!$ƶ��;�<��ُ�w����� ���]�� ڈ��4q�͚6h�?�h�o���GY�}���אtY7�Q�ȏC��Er?�O
���|�(g�����)�y��G�3��>������!�����i����P5�2FjN&dG=7T&xk�Ҽ���ߨ1�ľf?-L����>[O�h�9x�$u	+}�p)ӷ�j�"kq����`�t�7�C��(c.콿�1���m���_�Wy�n._��� M�&�w��>E�1������o���!�IX�2T9lӔ.y��1��vȆ��q���7?�됍�D9����\�Z\�C���=JqlF���d��3�"R�,�W��~��+"Ssb�~/�h!r�b��A�H��Y��E/z�}�����z9�����M�- K�9�e�O��WSZ��L�ʼ��ٻ<�"$�g�#-����/�[e���H�)jǢ�~��9꡵�3�Y�����|=ޘS}5�nV���~8�Y�DG�D'K�1u��oa��M����C�J��J2������Jo�n.��o��������L�E�h\��?�����ͤ�X�P+�o�6�o H���5U�o�yj"&�����I$lw-����r�Z\����~��Q1ŜFG5���[ۥxv�����B������v��z(& ��-��yR��7�Q*Q�w�i�#��f��`��r���󕥓��4°46��0\��ʃ+�IFsHX[�uaq1	�$ �W�I-~%�t�\�z� �����I*�,�b���f["�����~��{��4��"��,�ۛ��c��J�E���{*s��]��G��k(��&k������(���ŻA~��W�����i� o����1�Ӥ����4I�g�B����*�>��r�ۛ�Tu�$F�8<<2���{���j^ú�V��"��m� �8��Q�0�@z�0���,RJ��'��>���������L�|ٷ%B���a���c��..-�����-@��������
�aNH��*��aǷ�d5�g�E����?����Q}Q�D#ɛ�~ �m�tT����\1e�P��]�-'2���Կ0VH{�)u͒X���W�A�}f�O1N.������vrDs�+8�g�Y�S�w����5	��+d�՘Ч�|~�5?z@2�a\�f���ď����q�<���E �o/�׿y���ۺ�آqB��x�����w֙2�T�"%�#�]��k����H�1��i�kE���K�O��@�-Ѩ ډ�6G~9hzc��|�W{>�gT��ǃ�^"�I��XbDE��i����\�S�F�F~���o�>V�20�4�5��4�`9M+�7��f7�[}k�Œ�C��o��f�k?�?>U�D"��fM@^������oo�Y�ƙ�%�M�c��}�$�MQg;��|q�@��PV^Ϋw�K�T�d|�*����>D<a��������6�|���bdS�JK�^����jɅ�l'fBA]�銎.XM�3��u��|����PH����I�~���O�\��H_���>
Y������=��҉�勩�ExE��G�~�G��B��Qdz���T8g���*G��:R���N�m�rv�7b�\r9;��WL��
���e���=��aP��&����������7�Ap	���p�[�j_�O�}50FV)*[uio[D p�����S��aϵa�W�[�g��e�����Ǆ��\���,~�g��y{p�^�RmC�N`Տ��cKB���Dl+c�-�lzJ2_^����p���~.--mє��jo����ڸ-�HM%���,��X�Zk���/�Օ�Փ4��R��n�p�m湑����H����Lq���?e�BWU���m��R�)N7G�c)�����3F ��?��{>Pp�Û	5����F�.~�Sbj�N-���o	܇�Q7f�,j���Q��.p���zo���s��w�����Ԧ/�s����$�N�T��ԗ�X�Mj���fw�x�3���]��U_�*��\�M�{I�?��'x��&q���EJ�t�w�E�_�r�+��Q��K+n���tm!����"�@+�aF��l~�5M�;-�GGه���E�ѽ�۪$`���s&ఫ�y[��{��83���GK�rAAR��f���������9#]B�_/��x�oq.}�t���qqr�e\t���g;�~MM���V�qI}%}�"���MK_N�?��:���I�R���(D�%'�o����U��v���S���Ś��X)k����G��K��"d�a��H�:��s�V���H�$&f�n>���$�U9�c��1����?	�	�8��,7������no���ۋ�N�-�m��V�sz�v�����AV���݋��@�$=N}3�cI���P�G<��@#�V�����:.�޾[7�Ff�,�Y��_�G��oG�T,}u�z�W���"�^��H����'�r[5�oH�0w�1~B r����%V��c{�����*Z�  ��D���x�'7����T@�k��ѳ���~�=}�c��7���<A^o������ G��,��lUT�\^Y�=���jo$1�	mϊ(1%�	�Zl}]�|әab6�$S�*cB�/�ǝU6�dt�0�2�</9��i�����_�ۜs�o'�����ks�tll,�n(�j4����k~MA�)��ƀ�P�O�ݣ<Ή� �e��'g���:>m��em:�E�h�V��$�!�ӮD����O����w��O�R�,�i��m@�=���
��Ņu�4�Ä�ߤ�5U�<]/�A�$���;.�bc_�LԷ���`!�!pբs4���8J:hZ������;U9mX����7�T�_����7_���x�l+|L�5����x�G
���Ҳ��񋆊�>�tF�L��j����e\��D(0��~~��W��\^��>~wwwm�������7F�Y�|'�S5�H�F6�K���_�7G��&�N�'����\�&B�1�W�t���Cc�~�ͧB��͚�Ϟ=����h?`y�;g����+O
�X�p_A�,�)��9��m8\Bѥ�d�������Z�����^ĪҊ���Ú�%';;{�2���{۴�j|��m����m� ��헧�%N�����$�fA@F�j\�:<��*�)^�-��~�D/�L�o�Pqz��j�Vʡ�n2^�H�x��šV�<��#"�}�~HO��Ϗ+n�q��cN��_�C/��kW���9�\������U����!-�t���y���A�ʫ�z�p6V�� ���6�744�������dx���.T�,���ҨeM?�%�c�,N��C�~��6K�B�8�9�x\���n��qw�,X��m��,����mkW��
��o3��(��(((���2��Á2(jk�W��~x�090�0>K�y��A5�zU*����3��5�R��@ds��	naF�����6wz]���gu�J�Zr�����1
h�=�"��h7Un�����-�����4sss���d�}c�!!��~������4����^�q�Ag����O'�^�nGd�F?�q���^%���񣜍0,L���C�Ly��;w�W�F�GH��T%L����^җ	-����hj�<�W����{mX��ν��$;y{�ei4��w0�O�F1��2L�MS7�^L�$���7�ޒ�q.���?z��7N��&���������Ȏ��S}=Yv�Ug8�;-.
X�˗�C��.������ʬ@����g��@6��:ùb�T�
����$q.���>J6K���o���1���a���=��)	���*��|D�?9��Vִ��F4Ѵ�
"(��M�t���+�q?�5���'��F%�D��I�?v�����#���im�`���QI���3�D&L���$MW��j�����Q����F�1F�Y���_>#>��\I$.�B*p��k������Z����u4[T���ςW�A��2@�VƔ���I?~�z-ё?y���{�}.H�����{W��W_�|�UT%�������4C�K�T�#�5m��MU�U��=�󎰾
�uJ�?U�7U`քo�rr<r���%�v�五�Gk�����/��d�}~UPR�M��0`*�%/��w����[�/����i6�(����^A<M�ϔ����#�;C���%��*�?�Y�QN�|'��,V�k�
鎺��f�(a�������k�Hؖ|���g��X�������
>r�(O_:�.�H.�H��.�ۼՇ�pHhdm���]�l[j4�i�f�ѷ,e��<q���3+Q�Np�Wؘ�'�M4$�%��,M�)s�r=��X�^zQ;m�}��z��Wv#tC�]��Y�N��Yl-Ԟr�d�]�U^͟`B��P���0�<]Z��GxZ�� �&��UM�pܑ�{�)KAavU�.� }�{�����1�/�z�R�҅�d�K��9�)r�����*�i��]/����BY<��÷�<���f�b��tD������!�4'�!�֒57��098:���s}�x�\DW��<���$+�y�Cc�\��0hF���k~�c��x�<�� 4�R�W�9QgJ�%���h�2�.�յ�~h󧬝j/ݷ�,�Of�V�L���T,�ε:��1K�,��N��.֯k�#w7��~����{�S��,[��:�Γ��b�j��Ȅs�����a�f&����E���'�[�R_(�*h��6���Yf�)��it�����x���R��AY�1�M���"��j�I~�"D&����OM��mng�'r�"t����An��	��P�{����]�􏕕�I��WZh?}2�ӟb|o����>X���'���d)D���|&0�j,VAߟ�1������� )�D�����v��_��=6F�^)��� 6���ZB�R�7H��w���n!�.�J�$��φ.M����X9��C*�PЁ����m���n�1Ƈ�� |�3����CP=XS��*/�)�^k��<�QN^9����N�]uN��n�P+8@��](�]��F�n�Gj�_"ֳP2~�R���/h~��B&��ۋbX���fu���&&������-��?�9>1�3������8���j�1!��x|vZ�&~dx�[����(�>8 �8�}	4Q���� ּt7������:5x,�����p�lՋ��v�Z����PO񈗋��&�Dt������D*H�Q1�����>�'�LAV��'�l�+�!V[�x ��J�5}%T��H
`�)H���M3��9�L_}�j��V�1G$�F@?�������ʉ=�Ǭ��$�K�����vPN)����f:��ڮ�!�^��F�_=�
��H�K)>#�4nvn��"�S��p�h��|����%*�~���X�%j�]���Ӟ�
�V�?E�h����{���t�*��Fb  :��+�=mN/%'��
���I����ǿN���Y���N/�xO��M���������g� �21�RF���LڒMMM���ť�3�s6cc0b�M��	u���&ԗ�|j< ��G�H�!�t;�Z��k�2���^����۴����;���=|C�B(/����A�nG���G��Y	���3����2u�`S�pqVb�Xu��yh<:e~�&���%@��"\'ƣb�c���**+�"8677���v&J���t>�V4������X��1� )F���L��z�wA�ns�KDD�=��������x�RR!���D�	X����\]�Ҙ�K�'u9��;Ѧ�G=��*�1�9��թ�=�����!wdͼ��k6�9����!�`�2�2N/�*w�&��WZ����ɛɕQBB+
m=l��8L 0�j�B��K���K��)�1ch'��C�RTȤ�Z���xD���� ����"��x�FhW�B���T�Y��u C���ɮ����.�ގL�������RB�Au�]�M���+�/D�m��hZ�YS$耬�S�1��Y��2H�"_�@��9��a*7�!3���c4��R�M�r◇��prrv��)&����׏ے.�yn��]��2b�*J\��c@�@�N��Z+s/�a��_�Ь���d*�4.��9	��0h8���p�,塖ㅊ�����xD��w�&6�����S@M}�n�m���v�3l2"e'�����4��
�M7�ldZ�%���n=j���e�|�c/���
p@vi�Ȳn��r�zX��rR�E�jDx�����5�� ^���M�ej��o��(��Z��?��S�����`p�{��j�aԱ<��ν���0�����ӣAd��Dh?�z�$��l�����L����!N쌫oHhe;���%;���H�8`����Fm�UT���S{Ia��f"���K�=c�Z� �K+#2L��J�^�N[m_u��F��:�q�!<�:G���?+DA�a����O���L�=^���ܾ87��b5�̴=]� �^}<�Ug��p��q�p�w���K���Q^W������"!!a�A����c��hG�
ƔrЎ0�]oq��?"n�Oc�!�}��͉9 z# N��"�فlQިP���h��	#�j3m�	M��vl��fvS����QǊ�=+J���l���"�)��9Lv�;��e�օ&�]]]�{�����&J&v��|�-��O���iLP���ҐA5.�-ey?�<<gtv�1�n�Ú?������)FMC�2�
�����(qbb�z�R��
U^۪�E�;��1��u��[��;��yq%5;<���|�$1���b�($[�{6�&��;T4O�ӇK[��
�� e����%��򐬿�ty4��O�[��00���}��È�}O���b����ǇkS�7��Vhh���|ؓ��en�釃:H���0���NM&�)/ʴ�w�^��^��H���A@�x��^�W����;:�"��[��4e���Y�������+* �ezϫ��"r��a�!�O����%T��&��!��#�ɵ������:�����=���2x��h᪑d��˽`�d����~m�p[��p�s�32�1��x�5����^��_�!��;[|�dA�H��G��{1�#��Z4Z>��v$��t�\z�7��vr�\��'�������E�3Ob�Sl�sL��#fsV���Mk�ր���L�Ѐ��a��o2��އ�^���|#�x'�H���ch�a�����}��a�=b�����m�'b��H��<n�>s�ג� �$[�BU�uB�1�#�̶�ע��ڂײ�>�f�I6��u����	rV.�V!�������2�Y�`` ��a&�y��� ���1+j�2��8A@�����v��3�Ó?}��"�
��vw���@��<��[ȅ�F�P��%����0LO���))�Nl�h?=���;����?P�n(���z��@8&ʈ��bc��v���6��hp�-�Х]8��PYœ���c3jǾZ�����f����3:��d��B�l���ŤlP�6[y�&k�q:a�k��@�UqՂ.�fD] �~P�����cBD�[�J���TO�GR��M����J��OY?�+Un^��ed^^~��->���2W�{�����%L`��x����k'RԷk=�X	�&�A���ό��	}-�`��Yʝ{����� �X�p�Q���,�u�@ΉmȎ����"��]3Cj���e(:L�$�Vܦ`��FL�1������%���*�qK����Pc�_d���?M�Q��=��GO�-�r�8��4��<�7�*���Â��!_m���t�������[OO���`�c���aA}eo^T.��l�yM���i�燋�9
���~yK�g���_MG�~?���1�2��Pf�b������C����=��c��hM�d���G2V�H������e�$�V2n�'O�s 9���� ��k�����{�˭u(���O�5�:�J�I�3;� �C� ]3}�����0՘.E�)6k���h<B�/Ԝ�x$�Ђ�*\��"�/��`��8��H�a=cer�" ��./��W~�	�ct���
�W޶��m��Ca��pғ��]���/��"���$�.�p�_ﰦ�,�`N1�c0�K�f��`%3���>����Z�#pI"����]�M��	�j�;�V�p5e��$�����3����?�~�|����o4T��j4��2h�<�Q����!Ү5T
=|v?ec�Df ;��?���X�cь���l�������-G�"����B��.�K��"(�A�72&Ǌ�F[�g,ZA�E��JΘ������t��+�,T�P�4���I���K_sEOni��`�3ᝬ^jIa��MS�N���������,��#�e��ݩZJ;��xڟa@/8gs�;ß��ىz��j�������\M0)$ǡ8�'5�=�-Q뵣��!���)���l6���˂F��D Q��.O�h�Bn�(\�}�n�?8o�r�[e,rw�+��$	�a�4�F�՗$�]J^����O���4�a�ih	a��i)*
[�0�p���q���0�O:��8��-y�7D����3c4�P-vT׍�`zJ蟶��]j�[CL�JrZ��vHV����`���9ɕV^b��uh���ϴق���؍QO����ZT���x����ʠrI,�/�r���䜦��I}�/�[��U��!�w��Y�j,�s�Q���u�dyJ��I@��[��j�k.[�e��I~���I���^6�A�����{}�^h�\�����"j�%��>���M������i����5y!�B;���I��4��(`Lފ
}��6bƮ(cL k��S�ui׊���	�m���UI�냴�.i#1Zܿ���6�,�i+�)�:#�n���7�0|Z����0��~��d�F�����X��d0�����i틮��������}�uI��k���B@�! 8Ĵ�@�W�x��î�:]����(�|���/ꎎ;M\t�I��>�G�5����>]�Q��v��8��$9�Ht�_�A.�O~�m鮝�ӱ�)+��y
+/�� �TY7��D6����)ǁ�b�EPvխ��c}T�-�Y��6�Ձv¯�P.#lgW�Gh���jF8�$o�lM����/{����U��m��
^��NF�G�Y���Q�%�m9��� ;m���i|�\�����Y	af��v�(�9"a��M�Hy�£j�:�F�" �����)��%`	��(x�wً�C�����ȇ}VU��������\���9���7+C���V|>%�z����ٚxϥ�΃��#�8�l���2����)'F�#�]�O�ah��(�=�B�ݡ�?��ςM��˘7�E���D�yR��ǵf�C�.K���C^-į'�|�S^6�G 1E�U�8Ǭ�؍��8=wţ>%��&}N[��((�7�	&I*�EлP�y��������.��)�4��锬�� ;T�K�Q:�������u����1�+���5ֹ��<�=[�Z�X�=]�� X-�W��O	5��ţ�+d�K��?����5~����t�F��.TyL�¶�����E����׭�>Z������VZ��}�������Q+c3A�OG[�o��AZ�(�U��PLd�&fv�l)��["�~N���̟���^K�y�
8����;����th'wQ-S��q9�ns�1��Z�o���8����Ɵ,𿣚BaJ�Ȃ�~�l��S楆ѱ�¤�8$O��Z`���DPq(������s3��wt������\Ը�!���i�#'xY{�XQ���������	�BϞ=��J.@�6�B�d��>��u����d...�e3��8�wH������nV׍������?,GDn/Û��p$�a�{��9�*"��\qO��aL�(��ڶB�%<>%��������4���ù$Xz�u��E�{?%V��+�x\%��������?vt8��W�uu7��C����el�7�(�Z(���u%5��*rm嶉��>�<!��S�ݛ����W����E�����.g�֌�#Eq��Tfp�-IT�Q�5ޘ�ދ���'�.�>cL���D����\�u�[A /V�5��7�y�xI���\�Da�K��j��L
	���:dG>�ܡ��qҾa��vF=Cæ��u�Ww4q��>�%��qa_X5�p�/H�|����d&�B��%R��O{ӥ�u�|�	������'3�e��	�ʿ�YNÜ��|�zu��o1���g�"b��+Ym-C�q���I�vU����U�M(�����z"nv_9�WS�U�+�p}x����@�ŁQZ��Δ<����_�֍��hi�UӸ�ﰫ����Ǳtk��<�
bR_yp��Mr4������J����x>�����Z��H��^: �+�	�K/A6���/ޘF'�_�u�ڈ������4Î)m��{q�ϣI!mv�uv������+�	���ê{U�{u��-��J]y,:��gl�����蘘��&�_�Ü���8���++^k�M_�����	�����iq�˰������Hb�<d]f�a���w�ߑKBbfw����c�y*\'��EЏZsC���x���NE�V���x9��1��J6˵��Q&k�^^_2/��7�tjX�S� �Osw�ί�ǡ��T�v�'m}������Bu�Z����x����<
�D��ʏ���I�*XP\�#>��3���?�t�3��6�%֫XB"��e�c�e����N:��אu�E�*C���.�_^�	���N��d�,�	E#T�؀+��p0ٕ���8���m�N�S��P=�1p��׿n�/�f�|f�H
,Dñ��_����X�d�O`�k��ۉ= j|���u��ꄆ�~f�� Rx�VU�&�Y����.UR�)��c�_fӨcIx���W�&}^�o��0F^�� �9Y�3�1�_�A|�R�I�b��)7����%4��/��y�b�[G�/�a��G���|�QQ�x#�jD,لك����>���C���2|̩��-|�tM��23#����tsD��u���~8+lsӾxrǺ�¨���G��������!;��`d��G��'Dy��s݄�EO�׉w�.��nF�uR���4��$1��v�S�k�eӢO��xQ]�w��U����|y ������V�܆̯Z���)��VHg<�����gl��f�:䏗Gې;3��!�B���&[�Un㓃����\ܔ|�&;��E-L���
�irƞ�b=���Ox�t�]H=rRw��q"��퐭���b�I�,�=鉗y!s�Ҝ:ٸSv���m��a�-pY��e���B�E�� Jyu�����|&2+p^:�,�����sd��J�I��nXl�y
[�o��_ٻ�`�|O�����=�ܙ�MOO��'�I��
�0�R�|�aZ�w
�l��Ȧ��u�䶨m�)8	Gy�`˲��2ɭ�!��bL�P����V��D|�6�7�%7�QZ_{ܹ�ʗ�Qb�CS��C	7sڮ�Su�� 3M	%Z���N9o]�f2p�OV��b*���_W����.��p�X��$�x�C)�i�����Տ��u�+�4�*eU�26�a����tr�2�V̗����տ46v�3���uD���R ðpy��J�{�盐q��m�-�b
�e�I�
�$,p���n�eUQ�a[56D
?��=�8i۽����
 �'��xʵ����K�3�x��B,�>r�LR���)z����Ÿ}��u��͘� `|�Ƙ�����As�aԞ��$�vErW��pY󘏷%/��pۄLA��$�����я >(��~*Kaq�a�#���T����I����K��M������(�����Yb�ld1��,(����ޱ�# !��e������O[Av>>Z�a��)��*|/�b�ً�G��%�n.�<��v3H������0�'1��~�Y��|��A_����m��o�V+~v�|�C��T!8��/�C�tW3-���JG~ފP��$JY����6��_o�~��^U#���V<a7!]������r�1Q-��ֿ�����P�E�ܡ,6&� H��r�<8Z�y�Y�]�������"R���97�����˦N� |ӌ]�pD���l��O���if/y2E���P�Wg���U�����_6O�Q~�K�1���z�R}��!H��N��WkNK����.��&��X%���pi=�'깡�v���'PDv��w�,	�����WB��f���97��/Em-��~%JI-��{o�U%f!@��#Xo�4'��:�6�r�rG���ѥ���7��w��9����f��O*G�1�d���F5f�!@��d�����������ʗ�)d�d�x��]?��yz��.c߶����8��Y�t(���������m�~#K�o=0L�)�����ϖj�m�C�bt��1�yg�q|K�`C�~�=��ֿf��x;�q�Ld�����(��^J�H<�'�N�)PPNJ$�Jx�/'^v�v�K�=9� ��V99�:�K��8�����E�a7�-c��6��s�0ʢ�S�h����վUW3k�v���Yє& #�}�@�\��M�[�N��&v��L!Qkw/�G���J/�}g~&~n�s�FB��@kb��Y�\1�q��p������5s�獳#8��LEV��\Gk,��khHS�>aЬ��)`�=N�!��u���hekٱ0��Ֆ�1B(�t�ˁ#+�`�ځ�zN|��oN�%��EYcF��fL�OH��P�~ac�u|ϳ;1k]�����aZ�`R� �ֹp���*]�L�÷iDhU�����ҏ5kuTu�Y������$��(����p�����/l��
Ǭ=��U�O?@�J�h�y�I�����Ixr���~���Wo�mPQ�޴�������f���/݄��w*w���C��E�v��@�Y��y��]dv��T	(8� �72=�* B��R�}�����
�C2���㓖�O.���D�����S��9��5�;�����ӂ�zY�7������Ҧ-Ҷ�R�̊��������*�R�{��_cJB����}�y<0כ������`7_G���Nf�f�x�j����cJz�e��'�������]�#��E�ZH�I��~���h>m*Mdd�C��c�Ɋ��GH+��I��
=�T�g�0���$�]�bAY1�7";��9�9_��UT��?/
���$�7Zo�`t�V�w0"�{���u�EƔg�a6�C�G�8��YKxh4F���S�[�0�w�{���]�� �q�/��*�Ki%*����f �����j��Z@�8�t8��� ���BB��bf���@T�y3�\�'vS�FV	{A��a;�#�v��\h/Z��tQg�}z�jg,H���SC�����v��>��k檻(�E���B O��-������(��-t)�!�h]��|���j:v�VU��f��P�N��f�9QG��~SZ�n��K>q(ŢkSc.=���~T�c�``�.��t�Tq�&�^4/k�����l�\�e�'�������JG_�<��Hx�R�+��M��(9�1�ʢ�h���c�kP��#�o���'��4u
���M�X�������j�񂄲������L�4A8�R��y�#�������f��yo�r��^��>�5mbH�����=[����P1����o�;�(h(u��������K�Ə+�s޵1�,nCL��/��']B"�=�v�?�1��C�b����@��gܒ�U@@��:��L.y,�L
�X��Tpx��n(���ҧ���O:�Pmn���'�4A�2��I/ʫ䄞֮��	�H�N4ns�se��,N�C�6e�.�|1T2��`,���f{�;`��S��d�R���Q�ZH�����ݶF�E*s���A�4�Q��GPLn����Ybe��Ka�Ă�NR몡z��h"�sJD=A�A�M�0�^x:��:_;Ü{�9K_�Nio�fX���ZN����>�U����N�^3hu)�o]���7�'NnV2��>3\�z�r&�L2q߅~n.J��~�C��k�W�?�no�%`/��dˌ�~���5Pm*t�3�Bl�U#�u�*s>2x��l:J�f�`�x�U�2���Ϩ��$�e��$�E�jYoD�9�N/QJ[�I	���\�Vb�������G �k+��8��Fg��d��cA˄�b���L��Ã!�i�w.�>�U�Z���ؚ�Hua��͸��)ZbGB�l��|kJrY�8�dT�^�h�~;pu�vYJ�qm�0um��[���Sv���|4�W8�d��� �1�����{��4�t�:ϟ���a �TGc,E}fr�q�d��>n~�Ƞq�]��G��� ����̬ ��W`G�W�(\�.���$]P��M���;8\$�s�[�����p?�!Hpw������.���5[��U�5���ｚ�}�9΀�J}��
��g��ՙ=D�`�"��_U�q��3�wI��?HW��7�f.X��O���(�_d�L6�,��퓊�9t���o6�9��Yd��x�7�~��?����sI������6
�Ϻ?�D�,�8elO/�C}�a�N�k"�1�=�b����r$^�|X9�����1$� �eC�:��x�'DY=U_��KV�5�I�%d����������w_ �.�
ʱ�.B�TB>/��)M��c׬�:���Qd<=��w�����wLA�yE�2k=U�p���>���s��Y0Uھƫ�� n�{�H����X�$X���'���[�*����i��,��w#���I��T��O�Y�=�e3�pdl2��qA���(0{>u�\�+�"R8uw��YAw�5���Q����rk L�������+g��!�h�i��,�?|�Bv=�po3��`^��3�Cg�z�x����Q7m�����o_S�	i�5R����=A?N!�@������|�r�F4���q�&>��K�K��ی��=q�mz��E�?G6Y�K���<���!���ɫ�����Mz��r	+��y	)8-�eq_��_-Ƈ�ב�ˣe�E���UR�p�����3�N�Ǟ���
�#Cr�mb�RV����Ck�C�Cq5բ�'q ��ǎ���&�9�4���c����jmbw���&��8���Ԧ)��a�P��b�j>�h��%��Z��K���@��B׷��=��%7�oxy��P�K���><���e��A;ߚhd�6��v�Ụ1�pX�G<N����c����Q��G�bd�Z���C٤�$�&o�^B��͡jR0�]���8�\�3%A��f����R�v����_i�x��޲�_�D̡c����q��a}]q���N��1-�C/��Ă�A�߬ҹ8�댲+�lDѱ4]Ma�lDy:�1[<"R���ʳ�0�"���>;���S�M�D2�b�G���urie;���A�hz�%�6]Ө����h:�Ɏ���T�M͊I7�KM�O5Ywc��>+Z
D�;7mp��w�@�q����MTw�L&�'�WE^y��7��莒�F�v�����x0���J��f�+�!y(/U*	-�G�(��p�9a
�,>.�4��;�8�������~b��B03=�����Zz�=V1��?q3ʡ�af*CDv��a������Y���%�()����9Pe��x�ds��!�D����R���&x`|����FLՄ�o���F�r�~]�B4@�3Bǥ��O!)�����JAA|��tc��='Z.�?�*e_%�$
��g�k�˨33���*:X?� ����+L2B6��Ek.���?����0�`�1�-���w1��܆2�F�5�
��9D�����H�)��#2�$L��$��q��Z)����9+�ę�<�]ur�.↫X8M��>I��8�v���(���/ vLfׅkD
3�ă�0&�j|��-*m��ElL��/�Au�F�g�QC$�x�N���f!���F'*����?]�Kq��(�A⌥�`��jc�G�����0�G���-�@}(�/�^
��6ޏa@�?e��Л�E?�y�|����p��!�_e�=;6�i�q����l�� fI��g�h��?�E*�е�DX�F*R�Ka��jA2A	���^=�J�����Q�$��n)P�(%��d8��tj���� e�\J���
	�|�A�+$©@��7��:aJ9>�$F�"�������qa�z;V�#�LI�j��M�!_����L�Q�d�yp����9\�1�Z��j뵃�?AP�u#	���M/0�g�`B����a��:i%����Cw����e"�����J���A��xR9�Y�	`���/�q`�����ێ@{�gh�2��;㼨���v�v�O�P��(�NDlA�e3���9U��z���
����Ɉ�Uj�Z���; %���!{Z*�s��"���-w
�
� �6rk��T��%�Oh`�j���￼rm,����� �';T���U�ڙh-(06���~��r�)�`3j�_�@ 5>ٷ�V@N^�Rc�o	'�i{��8Z-y^��ĀAP�{Ǆ�$C���ٓH9�HR�Y�4m��EQކH�����S��}8%<K~E(M�F���&f���2�`)����������<��Qf͋��̏sN�1;��Z�o,�K���Ⱦ�5�g��m�#����d̊�\q�Iчr�s4;W�/�V�U�i��t�V/��³�Z���f_q�G���_*��ś	��Q��#T��bE�ώ�(w��C��t�(Z1]~.^���L}�9�"�a/���/�Q�����W��W�Vs��	D�cm�f���I������͌r�3� jI��fO�t����*h|��8PN��˿)���#x�'��w�3{��<�l�Mk��s�\�b��b�r�Y}Y��yiޭ���vSi�|(�� ��cE�4��%�
�'� >�2#�{��9&R�����#iZ/n$���E)~A�[�!f#�+�ԂW�6�+';|�;�YP���O x�(�}���"ώ
����U��V'##�,����Z,�4FV��3:��@� m�ݏ�y.�т�vN��gVc�0�0,Jc�~��rCҙ�p<3�����6��H���ΨU�g8��T������?�d�a0ؔ��_����$�)
e�o�j�Cҕ��FgC{]�c:*�nCdDQ ����)�Q)Vj6?YpO���խ�q�t�	=ַ���Y�5�P�Hnf���q�X5c�C!F��DTb�6~mK���x�.��`Q�����+�8[7*7*&�� 
h�韡
Ǭb�(�믚������׸�K���,�]���[5&�BJ��*'� �S���,�EƘ�2���������б�������U����;7�R�AP� ����Z�(r�����X��,�R���o�e=�/6DءI{J���g+�ð)��x	7�h�WQmf$~�,�/��&B�g��D�N%:�6� ʟ�Y;�C�+� S�R����b�H�Ã�<�9�sN؉��4n��!�`�8�HPn mؽt�]�T���_sR.27�/��ˡHaQ��R�$jv�y�Q����(��(�8��F�k���VE�V��v?��`M��W���3TN9� �0�)�p| 
���]'5�dc��q{k�C_�S,�߄R�� �-/�I��/�͝[��p�A�c�$\�����0A<(�W}'cx�t�m����o_^�xv">��X��w8 ,7�ԅ�A�M�������N��k���bOZ��t5F�Q��%�6HL#��4��

�Y�Ei@�q�K���w��K��H�h�Jb(Y�L���Yv���jr��'�w�$��*$<~$��&P�?��%�FH�1�A��)x�jQ�=Rp���chՊD[	�J�T��t+wU��k�˷��q
]�}ؓzWը�/-pRu�!f$����6�6͝'(@S�k(��c���C�c�CEDz�I(e%+	:`ybbT�﬚�����A������>�::ΔMЅ�Gm"�߫�����iٗ)s��S4���u�ĕ'ǫؘ���Ǝ��0��JW��c"�,$�b\�ĥ�H���SB%��9�O��.齜�~�}n�K'�o{X�V:��n*t������NBJ��wl��&���x�LUH5���Ȉ�7]����N޿h7Ҷr�l�{x�M�^/��L@_:�z:$g(0����`�X�q緩_����:JD�r?g7T?g*��ɼ#�ė�͐B}��Op�Ã��߅�G�46feV�x�p��$_4]vDH����w�s�Wh��o����f��0��D"�l?���E�!\�Y��~v^���8�D��a.T��{����!���{���*��������D�s��8"�oӫLϑ��~ױ�xʬ��7���T�μ�gbp��P�$@�b'��DDԐr?���O����,(��"r�$N�%X��s�����EI�G�E1͔�V|������w��!nr�3�%D��mr���?mb�=Qyn�R�)C{(+�b&��t�.V�b��-�ߘ?���,���Uz���oFA*�o�qP�+�0-/�A~Z|��Š8�~}��9�ܪ8<��e8,�*�uiGN"��1<�0�����%雳�WG�U:���)7�4��d�����aJ.#���v��Rl�"FM�`76~i۽=�റ��>�Q������g��]�����F�J|<�l�X�Y���{���b���+w�~C�O��Ɠ�f:���N���a�"���Xr�i�2�l�����{%�J�������Ĩ�ZD�}b���7ۉr7�f
LC%����&�ʼ4y�LB��Ї*)�#\ڮ�ƞ,�"1�iB��n6ޘ�����d��u�Sg�G�8�@nG���$M�H�|���l3�''��s�m�Tx�C=#�)(��>?�GsΧK�֐U*�c��|N�nn����RțYr`�a<��޳+�0[*��%>���h��4�L%�(�E��qݢ�Qz�.B$��V�+B�8�SIsS ^BorQs���Ӻ6�t�oWo�,_ئk�5�u�W ک%��޶/4{����k����EC��\��������\�U��#�2
�ɵ����o�8��h����b�y,�C�1h��4^*"1��kc<ΤT:�&��[�wB�;�>��D&�j�x���E��8%�XB
�C�J���J�8�IV?��!�E��ZOi�VZ�i\��� ��X���>����\��)a���.ȹ˛�p�
P�U�awo���+��U�\����j���Ot!�О��p�L��_��PE��M�e'�լ��u*H�T��s�r�K����Mc���-���d�a��Ŗ��:)�T	 E%�O��w�
0 �a�P���W�]<�N��̅���	���pB*ϥ��+��0�9?��E�^��7-2�Ź�ʾ{��Ћ���ٛ�{��S�C�,�����|���L��6
��,&��RSܙ���H�/G,�Q��=��M3Ć����Iq� B�~��,���k�I�����n��AkZ��5B��Y>��Ɲx/�X�E]���^N�6��������|�tB$��au�E��\(�l��3.e���t�}i"Y�׶G�x�/��.�s��5@%��oڅ%$ձR��߭y���z!c!�-0���'ˋ�	+���:���o�<�)�xv/�8�9D	��G'�?L֠GJ���{>_�(���ŵ��s�=���7���m��+��"��+�g�|)
�^�J�_�u���&�R?B�3�z�,���Z����XK�,�"�םa�kR��8��إTDv=��q#�i�?�{��i�J�h���n�_���G�D$^V�պ���X���(+��z'F�iu젭�'d�
�%�M�UD
DQ��&MI��i1�.�k�"=��"+}K.���y�ϻ��iL<�T��Kt���������|�A ��xX�I�U���it����0�Ǖ��;��uml;Ȉp{��/+"�d�͞c5��@�ȕ�{�y��H���tV�5&$���S�5�!?�ݰ��ò�
�P%o�g�:�7#���̓�����H�2��1�Uܪu>~;y˫�޳���/v�rۿ�Y���yIMLL���y^ĕ��6��Y��ި�0*����g��F�YI@I����e)�x�"GEiy�l�Yd�o!�ĆP�]�ާ�iʊ��t�NT�����{	�����A���A�����-]4�FS�"`����g[�1#�ے�98 �q�q�}�����c�zцV�|�2�_)gBk95il�Ue�oP���^8�v�Y�T\�FO�l}���v(θTMH����;kJa.LW-�u�.\��J�q����^�����-r���_D�5���Yh����%M�6�\b�`�u��X�f���=|h��n�$�u���s�4z��ns��:[7Z��\	����/��!ai�4�@X�S�h_��M�]��'$:�?=���)��Ұhc,x��ͳ��1��� ��s.]�l�ݒ)���1�
m6_�J�4T��`շ7��WJX�N|Ε��C���&��I�l����#��1nÿ):�)e��"'+0��j������k�j���n�q�>�,g�;�cl[������m��=��UV��J�gޘ��jKH8�(�뿾f����O$�$y�q��Wx�����YQ�~�r5HN����7�-�99>(��e��Ч;��W�$d_gH4����7_��2�_����cfs�Z��\ֱ���p�ڄ�+p�"�
!�n>1z�*�#8cWOk��.��W���^�fE{����ߴ.	�������YF��pe�?HmE�N�Yv������ӎ�����p?�̼�z���/�>g�ߞh�;�>S�F�]�'���FK�2s-w�6��F��2��ws
b,o�W�ʫD���:�7�N��>�9���ctP)���SVwb�KTc�S��+�ϨMǃE�v��'aN��0�+���z���E�#��3�j �T�e]�q���q�z�=�T�ʎ�еlǠ����ɨ���=Ph܍�ڻ���u����r�A�5õ2Z�slx�<���(_
sւ7#����D��f������ZėY�st,������4(��I}B��G�n�v��(�ǺT5������|$�hӂ$jT.Կ3�6��[�-4V���������#C�вi�il�9�DXy! w׵�����?l��+����uBH���#�������D���L� dވ����T��.>">�-��C$�p�u�lᔈ����y�����!ƬV5�À�b�.M��r`y]6��`/�����]�2���:�׭���`Mꖄ��N�����+�D⑪ČT�c�W&��+դ923�}�~��?��F�򃬪ui�t��BZ�/ox:���B�M���s�Ѽ$~�1�*�X��'����ǲ��D�.�@��y��-Z#�s?,	,���z&i�|�3��i��G�]�L���O��-���)� C�p5/H��Ā�l.���{�.�Dk]�Q�)z�>"����o��!E-�j��2��Hv5����N�Os<b��_Ŀ9�[���743��Ҙ+�^O���#���,�>��V���~d�Y_L߈��i�$�}zfδ��!�}D�\jg8Xa��a��׶G�P
�/)q��#Cr�Ž@O�Ϡ�W͟6+�4�����Q�6x�մ��	��w�Qa#��[^�X���X�.��B��!8��MЦ�D�0"��n�;�x��U͐8�}��"� 1Jy�lJ�w]n}�q�p\Ue���*(V�c�=��J	����N��k�x��,%� ��?���h���&]c��>$$�i؟!�q�ә�~�{�)�p��8^`�s�����sѫʷv҄�χ.�Q�QE ��t��+�4�fv�Kg=N�Q �r�e�%�x��Ax��fǵ�|5EYݥ� ��
��j,����ı�";�.;H�MH~��̉q	��1;j̉���cn��@�΍�;E�$�O��V�jk��x��y<�W�7�KP"*�媡�B����f�MW��q4�i�E!��i�3�QR#8��p&�wOZ��g�mh�U!�t���{w��$�)��=�O��?7T��"І�����u�̄}ߩ�
�}���ۦ`�#4X�/��X(��XoEd���i\s�z(_�~%�������]�u����-�_�oNQ`Ɓ@��ܥF�f�.�SCHT�3V,�RÛ�7Wj�'1�H���
|�No?(�G�>�"��x��q�X���\�*5�i��B�Rm���
��χY�XI0������Z�J	d���\K���鲳?Ԑ��ɹ��6�l�{�p��ֺ��)}�V㟼bn�]�a�n�B��Y�P����w>�⒟����c8��}���ר�g� Ŵ2�,��{�o迥�%X�ء�� z|�$��f���l����xδB���<�\��j�R5����.�8t��*�Q<��Rr̠�z�6�Â��V i�h/�ވY�LQ_����(%td�ZY&֘x���V�gw�m�g���k�]���{�'.7����jX򫶶�\o�?�����*�'p�+�1]c��;���+�{WCG�'U8�3�0426*(�.��~9!��JT�8�ф�̏J��k8ӛ��-��5��H'�}�k&���*A:y߄ɑ#4b��N]�4!�f|E<� ,S�)ϩ�z�TM��)��I"��W�B��m_��+�օ[�&���x�������R�s�.����w��l��%~�a������	-��c}����I�Id�}�,R��%��
�U�K$�ce5�.�;er�MƎ��q��b�\[a_�,�C9�{(2V�9�������������ak��p�
�@����`!������r�� O2�,#�����M�uY���;|߹�ҽ�p��f�9j���h��|w�W]����}׿�����%�5��՚��㈶���j��5��0F�>	��˿��w�$Zp����]�3������F�अ+��~F�v��KG���HCJ��K����̤�س�&��ǹ-����B H'�O*T�u�q��M��%ޕ�ULs��1�ţ���$�1����M���|rQ������3���V8�ھG����;X�v?���3���).X��)�/�)%d�T�E���Bc�i����j�~
	`����}���i%̄��o�(ٴԊ�[ą7:��1q�~�@	p�a��:�Pl��1�d�OV$ʩ�L������6��!Q��T�|����8G�k��k!����\?��ES�(�xv���O�"�k��	[�4NՅ���%%�))"(]�*���lE�d���=Bdif��b���S���k�"�+���u��2$!P�1��[�b��:k�-�,���W[yV���t�̂J�xUb�Eх���c�$*�>��+f�l�^�1�1�?]^r|��/��H3 �&g���!,�~�ZQ�Ȧ�{E��Ѭ�e�ծ OV����M~w�z��g��8�D�TT�z�x���f"�<��T�$3$"J��_!w������Bܼ�RU�!E�a/�E?��M>.����.H��&�� ӌ�� uD`t��=Y &�B���,
ZHi(��2Z��{0�
E,Z*ѩZU�著��@������ħ3 f	�Z�5t�"@X�c�?m�Kf��m�황�{��x�P�����mcA��TV3�.�B��&��%6BY��TՖ��9�ϗ�	M�|����w�_��@�y��A��@*b����+��215-4�,�K0�/�q���kM��Ƈ�c�5]ڏ���n�ATf���\S~��"a��\1}hV�`o�%�sD�����H9�@��2L ��fV�P�#ga`���T�,>�Z�O9ZV3��o��¿�B����NƘ�V8��Z���Z��'��C�¯�{#P�?��[F(��7�b�镝c�?྿��A��Ys4r�~mz����р�Ti����ǇN������<h9qnK�*�E�&����Վ�w�"^(�������J��M��`%��(%&�ƻ�M�vQ�ƅ�����x�n�%��_�Xy���&k�=�%J��f����4jP&R�b�� �@0̘��u��n�Fu�ey�OQf\��.��B�Ȍ�I�,�X� � �Y6"��+"�z�P�T�w5����F�jث��.ЀK'n)��X�z�l:K���ׂ��4_/X�����H���x�aII>�ȟO5�>a�/��\o�A'��}xx�^�~<33���#�L*/ �8|�W�1�{�8�B��f�����I�O^��ۼh7ҕ_�d���6x��;?^��>B�}Ojl~���P{V�Wt`m,�WƿQn��i�@cn�|n��WQy�m)U$�9�뇙0J��V���8$r�4yxl��犚D ����U筄�A6�;;ޅDW�+�)d�P�Z]'v�Tl�p,�7�� �#ʻB�^����ST��ﴯLV�]���X��u�f^6��s�E㣣����E��L�j!�pq�$\N�">[���z����JQ-��e���I�6l<A|;*+�b�D��#��_^��#�Uq��yۜ�M`���z"&��	���^W<[�?�c�+½?�\~��g���Q���d"23�54���.m���;w�BO��[����bL�m�AhNVAp}*��ZVDݰ?�ܳ��"nFQԺ���Kj?B�=�?�����`f�j��>�c�z@EV#gXn'џ�J�8�xc��Z3ϩW�O}fI;��c��f���# N|ڎ��3�u�jOT�K�$Z��1�!���zQ�<��n|�eO�0d�z�
���yBn�'i<vX��,l:�%�K���"x�j�r�<��9��L�K�zѼ�H�:GSa`�(.AH���r!J��ia��r��]��J��ЌYE�vi�<.|z$�:��T��9n8_�~��zؒ�w9�\��W��(���Z��mXh׶YwȺ��8�x<��P񜨷�4��"�./�
?5O�o��D�!�� ���l�](V�prr:�g"M�W�*̅����3��	���u�n�,�:Q�!9bo7�_3/�Jte	�,'ט����8�Y�aX�+O��Z�]en�2=����|����c�Del�W��br����PR���W�����J��(��BJ�dG�	�	1��nLX.Ww����X�v-�P2��9ح0ݾ�����>�Ho�Y�0=�W9n���2��l!0�+�6�Q�a��F�J�$�P@�GG��F�J����8�
���$��^s�"%�B�YM�/iG��r�C�f&Sh7�ENh4Kd�Q�ǔ�^"�:���V�����H8Р\��y "-���W���	�s|�1�!Br"Ģ�2��R����~Ҿ�p�z��sz����
�-���I�1�=���r�uQp�=
��W^�2�vk�H2.%���U0ML���WH܄2�N�H33���}Q�Ɲ�x�����0��&[�/�(-�ӕ���	62��I9�:������p�IY~�^�
RǛ�{Y�%7�e�\y@zB����3�aɇ��OJ*}� �X@~��̀�Vri1�uͥ����}��1`��}T'�\���5MLv�N�׷�#*GI�I成�� �78jP��	�q�˲�'�áa0���K9���0�%���>kYtQ��K�t�(�/*k���P!�2j�;/��/)�O����ď�i
W���N�H4?��!��4UƩ�����b<9B�/1 ��b$y){4��&���f�0`���T�kv�S剚�f�,I��G����+$�6wO1,� q�x��h�u��2r�P�S������Z��Θ��\�x�Œ����Y�o��_V'�ۥ��='�|�m�P�8�S^��Z�v� W6e�fs]j�w�1	���*L����M�sfϓ5_�{���� ��������Y�c^�5���F㛙�+���3i�j�nuV.��������x�Ij�8.�('4�{|]\�s"s��em~||�����L�f~���M\�Q�9�����4	�ś���/�nm&0~ks�6����K���+�\ê��+�B!�nd7�/�~���Ns��y$�?�:/97��#*�^;�Fh�<
�/h��rD�,+�A��M� �v��_P�SOle�*���ک���]�|q]��<�-��}�{4q�!��L[���F�L���5�	����<<o����>���N�e@��N��~�WF��|.Y�"�HK	��n\A�U\�M�[��N[ۛg��6!w*��B����M���.���mnq'��|��_d]Ȧ���w�s>����(�>�z�f�j2a}��!|���P[ʕk�\,2	�a�'�hq�1=Εׯɴ��_��B��Y#�ӷ��Q�B�w���'��j����.���{�������춵jR8�h�>���$�'<y��g;��,�?B1���H9�b�g�����y��F�rC��K�{"�6�޺�f�a\�m��_�j^�x�#��4M���eY�K��E��
�f�L g2�a����J C�缤j���Vo�l܆X?Z�0��-�W��^V�n\wRW_O�8�o:�_��U��=�)-f?�bSFy<\��R'��6�g�=��Q��ʺphP+��$UZ���@��=9�������(��M��v�r�fi�S��%��QL)iօq�\�G�_�>�U6��'ġ�NR(�cZ��WBRss��
��N���2�������3��5-��� /^���y2�%NZ&N`D!����PL��#.�Ƈ���bۖ5邝ì�����X���cN���M���!�t��0s�\���yE��3?Ѻ�ai���F���������O�)Vie�3"�R��cu�9 `<X ���L���8q�8}��ࠎ��pd'������Q�Y��͔�
��ش��l9i��B"L��h�n{��1�ۃ� �1�Ls���^�C3�N��۴TꬿVGqD���Eg�cMH�H��F�4��R�o�~�o{���z������^5j?	V������p��=��lgV�F���ɵ+�Q��SO
ݒ�c��I݄y��>}k._q�=M���sȒ��(D݆n�x+ �3�'�@�3�����SX�ȏQ�4�5�w��=>-��X�sZ7W��
��ӄ��OEfWV�LN���������F�'J�}.ZAWPN&�kWr.v��ݢ��u��x��OV��t@6x��ճ{��`�~].��J�}���fZ&�*�	�-H�"�� J�����≋��.piz�n2�&�x5N�W]	#0Tq�����,��IوRp).�c�tB&��Ô⋐�s)N��!��Kxd|�H�e������=����Q˃B�RM��I�b����~������b�D�b,��=�d�d+�f-Y�<_�b��q�2��4y�~E*R�}���"�y�3�y*�uMgF��浵��Z�"��("�0�aW��XT\����X�bQ\��W2�e��Wל�DJ�1��s�:����I+�P. P!e����"�����V67G���0Q�m�K0��X���$�S�|��$�W��L�A�#����G���$� Q/�Q�GSS1��WUy�:3��;�	ޮf�m��q`5u��/�L���&�B��̇(��#T�ǋ����WXM�M��� a]h���̡�|d K!�NM��󆽌���+�M���T����!���m����K�U���ѱ����GÎ�񗤋sB��$�C�1����쌲����Ob��t�D]ݖ}�]-��������*�%h��ꦅ�6���h�L�&Nyɢ0~Q�V٨�omBe���������ڞԊ�
��ֿ������-����t����uD��M���a�a��RC�lP���*[8O�.��"oqp�6V�2^e���pȚ{|dt&o���9��tǙy�3|Wb������}٢�C޶��i�¶z�]��B�x.`�-�ѿ��F�e+�����ߨe1x���:��b��@�-k�ti(W
��~/P�N#�5��� ���������M�Ey�gE\����J^���:+�H�ߥiTy��#t�Zщ/�S�}�Pj0���`� �O��M�~�q�F*�+�ǳ{bl�$��Ev��NF���f���[7��O�MsO�d��?��Y�����R� �[�`ˌg=���X�=�yY��HrZ�C)т��&}+�-�n��C���g��~�rT8����N{/������K��C�����\S�{�����`��~,11�|"�H��g�p���@�;hO#�X��$�j�s�dտ8b�p��}l߹{�~!tn��Ȝ����	�� ��\�W��x��DH&um��4mm�FM�ҸF�ʙ��I�V���ߝ�ws�p���Ca�P.�j��]�o%|t�(��8"C�J4�ads�k�?zcOh�k:�b"Q�2���C��6;r�4�~)���jO��iɔ��U��ǀ��:G���y����r��C����q=��;.��xWfK><44t�'F~O5�RjS�@�N;���ُ�7�%��W��Nնi�./1�$��ڦB�fd"������J��I
'�Y�q��|��"	o
���<���{*&�y$u ;�d2�l�X�'�{.v?��h'�4�{߼h'g�������.f�m���L��|�x`ΐ~Hy�=���w�����J��DA_�x�?���l���VՃgR�9�`m�ʔ0`v3��!�\��ݱq��Q�X��"v,�߬��zqV&��Q@��h��͗g����>�?~x$��]���Dv�cӞ�����vs�#x���ө��g�룥`��8Y�u�p�0[�
��-��W
Y�׉�=�m�gn��T��)����㘆W���5|cU���mV��vk.�ɝ+��<2.iϘ�nf��q�鐓��jK�]�|c>�S�*����$o=�{\��	X},��v�~1�z�;��?k�NGy��ȱE�V�@��z�cE2�=���TI�Z�Q{]P<�p�)�i�����dȨ��4��nҾ��	@�_�TKu�^�C)�]�S�o7臹݇v&1���?}/z��݌^���xMuw7�lol�
	GG�v�
e�_�t%��(ϽM����;���oT@�!��	�������M�bPW�Ͼ� �	Pﳭ��,&\��%2T{�L�'��2�_!xN���PkoP9j ?�����i�+����[���5+k:b����gNK9v�K�@�gdL9�9齛v;�N��m������%��t�¨<�*��AI���
������AL��P�n��)�Ў��O��u��`"`X��`N�~�i��Z ��e�������P8���4�)'���9е�E��v_��444�9t�����Z87�YA��O)Ѐ~��_���l��C�Vk��bc�n�.��>y�Z<\����K�r��%ƘX�b�#�?eV����P�Ն��k�p�Y�-�62t������2�j�~瓥��
n�[�߿�;���[�q�CqYq��Yƚ�?�J�ɀ� :�M��E��r���@�:<��dEmkC`����_�9����R˫��ΰ��*�����k�˅�P��QV�K��PS��
��(����=(E�GLჯ�$���#�5/�r�w�mNP���4#��(M�:�n�8��g �D��3���ԮQ�Уl.�e̦q�co/
1}[!�
/�>�L����P&����\�����z �v��Gӡ5f����:���?eQ�h��z��P�;=$��"�Kj�5ؐ;\�%k��U��������N��R$��_c)+���)ۯ�[�џ�8��&����Rfך�\@#����*�w�X�6�֖��fQ
JP�A ���H���
��4̂A��"2K59m_�*Ae��B�+�����;�p8Xb �=��\�_�W{E���-w��L%��	���[�Tz#1 �䍐��;?[=��p�6U�ӫ'@:�B88 w�1`:5�^��Գ����J޸��z��T��T�fqH��AͿ<B��x���T)?`�d�a�NX����.�ԃ׬�J�)*�V�u. ��d&x۵_A�2��u��xn�](s�"��b���afD5�f�#�s,��J}�P�LϿޞ6a��u�";�h��M-��{��O�����)��������9Rky��\u�������e!a��~�"H=q�c��m�j��<�Uس&�N|��[��A�����?��g"o�Hogy�mV���[[G
��̃����$��9����$�`���?�L�ˮt
A�8���]~T�R���#ɟWB��m��i�"m�d���Xn�I�7�h��@1e�-_u����	?Yn��b=3�o�O���{�u����T�&�M�qJ]��e.��"yEב����ޡ'�h7I��=y�R�z$nʐ���򜣨�؜1U���,��	m!������x(�>k����<�V�ȷ�E(Ct���l֍"����W���[�Xq�z�>`1��r7�v���dBU�,��2U	bo�n|tB��>s��v�
F�R��z�p�<�5�u��T���F9�Z�r������Ȉm���,��λ�h�4��x3���0�j�;���0�������
d��Q,��W�[GE�}�À���� ��
C�HI��4H� �C�4JIw7(-�"!Hw�3�?���]�֬uc�s�~�8��׏G7I��>[�z�y�#�zf������T�:A�w�`�S8c7x��jK4�$x�
!�}6�h�I���
�穳�}�ͱ^Y�� }	(Hc�d7�A��� �&9:��洘�K�Ptj�D�Ίx����*�JT�\f��7��h1F���E�9�i����P ��=�o� ��AP7u��"8b�Mlޗ������\�ff��k�3�rq>YÒ��'�s>D�����>�z[[�*��D��v�1r�.�*����[&��6���4����(�V�zX�U�#l}���;�^�-�!��x�G����~C6D����[���j���������������ڗ��"�
V⫗UG�s�u7��'�ʺ�qmM�7�Ġ�[�G}C tJ���Gڻ��L�[2
R\1��9�",y��~����uM?~�E���=ߑ.auO�X�_���Q]��f��~V���L�8�Ji`�o �����Ԗ�yW�x�$y#�wD� \�:�]ߪ��~�A<JF��t���֚}�O�;��f���&y_���r��G\����q-~G@��df�rd}�����z�p��8w:`L����
KrqSr��C)��}Ԡ��A]v�oN�el`�����o��V����x���Qĳ���0I�r�Y���%It�eJǯnZ��b���#ԩj�yw�;��������Mx���-}�3�2�����&n�{�h�rc��?����8I��E��j>\0�~�ڴs��I��6�z>������x+5EffJlj�9��<>N1��Oۖ�cbg�]�뻢O~q�}$�4���`�AJE[���zqs�s�j�]�	|���XA�p�p���Ś%g
rRa�q��qJ�UmS���?k�'G'��A�P�i���}w�_�z���u�>�x�ґ�EX����x3��������Z�8�_Hs쌠v���U$����-��eV�=�<�@�v�lLL�1��Z�����sŃ���pv�z��n�uDNW!'$���g=t�[��lÆ�)�ݕG�b[PF�0%�Q�qZ��tl_�9!��0Q�c$������\/�r�f���V����w�pG7���c$�^y�2 �����ܟ%N����7?�S��s>��^)tl���$d�SVhS�;�Q}s�O�9sǺ��:^�w[�ضY��9���-��1�E1�A�Df���Z���ر.Ϙ�)9f�����nSœm�.�(D�U�cfȸ��iz,w�\�e�%ξw���\3^�o�+>.�C�
B��.�ZDb��R�/uw�:ϳҚ4ѢZ�e��|����\a�g1�5
�g<���[ȥ�,/5:#R����xO'�C����y��r�Ǧz?X�����q����x��9w����O�oP����� lJ�Us�4�*J���)�8�=���E�Z����Y&�йm4����pso��k�GH�?�/{���"�Ql�z�o�� AZ��4y	=�p�tʠ�D�|1�,7/�dA���aEb;�xb�}T��E(��p���oχ�� �}},U���)�+&٦���w��a[[V�M��~��<��������D��w�ђ�5������:&]���K��=.�Jߎ�]Li�E��A,�J�$g�q:숛�K^���B�N{�\���Y��ꝙ���/>�#�ʪ�Z=�J��VŔ�n��T!��}~�I+�݊��R����x�![[�=R(�nȱ����B+R}%۹�qeaYl���]�g;�s奋��.���S��o/>^�L�2ɃnF�P�YU􋊸t$�{�"Q[�~�*D�4d���؊�)k>���`�4��i�i̡hB`�!n�������pY���w��Mau���uq�k�d�&�4�͒B�Ԉ�RbFT�#c���%V�L����5 ?%>m�� �(|(����c��� ���\����5���褄c�F�ɭ���)����555��8з`��m�zoX�&B���O��i)�T��FjC#�]�޴�"�֞���r�Ο�+��]��},Q�:�� ����%�n�|ҙ���ws��
����ee�ZڡD��o���!�������xh�EU}!�0�/�^^)ʯ�U�5�p]����6lT]�5���ul��܄��4�
�b�!�ֲl4S�B'���;*��$�
�#��'U:�%*��`#C��r�@�-fIY5B0��@0z��!T/|�F/���)��mm�՞���+U45;�nQ�BK�A������=.븖�@ף�pͨ�� �|�?p����.�{TXe��8Z�i@�<�I/A
Z%<���.���=�t��?SþFD��'c���sMa!	-�c�@��C��fc"�P���ܵ�TqB�Xt��eXf=��W�t��T�_�l5a@���i���}��'�o0k�(sv c$�/޼e��9�����|���V8�lŠ�~0��;�%�T�X�2�H�EVdd3������� ��	�`�}�RO�xZ���
RNd��� V����?b��#tWl����4��aS�'ޘ%H}��T(��Ċ�U�)*���5����wA��D�JXoH�S~d7�=�N���U����ղ2�ܲ$\���������h�ݯhͪ9�y���az|'.!9�$1My��e����U�W����H�!�N��]T�,^�K-�FU����^�0�V�l���}d*Y�r�'"�����tW�j]-�����3S$�Ub��q�egog��G��Q@4'�?Y�.|�OTt�h'�7�a���HB\{vm��sr��"~���>�	�qr�A'���S�������.E�ف
N��˵���7���X~���ڝ�W�:{�rϒ��ֹ~�0"�Mz7�<$�Zî:���1vN���'s'{��T��6�����^�kɇ]s�ٿLIm�S5a�>�vU-o+��u��5�
�G1v�ֺ����:�=�7;O��nM�L��u��
"!y|��hק;�<�^��7?s���כ�]k+�M�<Ϋ����e&Q�a�B��<��Gw�~[�&?�rn^�	ɣ����0���'�H�֘n)^]M�խ/i�s{�:�F�>�y�Z����n��Z�� �G��/OG��^t�I���=Tz_^��W�z��2J�t������B�v��+ɳ#z�,�����E�!��(�)�J��R�v��/a��Z������E�`�S(�}N�"���¨w��ehm6��]"qi��u�-���Hy/$U��.����zl����]+"���=ݫ�|'Q�n�C�yc`_2�έ��d�w�V/}[ܠIsxY�����%��n`{���F;���9k��ld<*��o��DG��|��e�X�&�H����[`��C�Q ���1|�h#t<�;Z���fe��,ׅ|�����A�4��e�4D�t�[��^z�W|;������/���dr͂j��S���k�c�ѣ^�Pf�/b��Z����$����ɧ�c}L�a���^ߵ7�ƽf��G}�~V`Ѩݜ��5��
F�_��8��|6���琿"���e�Ŷ$>��_^§}��#��q[L�at}��{O���6ޣ���Wȫ[H<ܳ}����F2;�g�J'2@�mc��v��;�X�<�f��2`�WՎa�A���(f�sadr����SR�M$�I.y����	����x��;�5ЛR���[�.����٣��Ǭ�;�q����ߎ��C`�c8����=Ÿ�ƴל�c���2�魣ɩ����������W>�iX�jZ1����i�,���r�Y��'v�<Lsۣ�\�ԁy��?hy�J�����;�D����H
 �F�ia�)�#��*��yu)E�J�C�\�1��5����]��fh�|�D��<�zI�(��"*���-����'�j�O@U5+ͱ9�1��1#l�}��:�;~7�ڂ�J��D���r�'�Q�l��x<��--�0�ρ~�d�5V����7%�s�w�/	T�r��c
rڞ��_)���5]�=*N���֢�qf�ߛsk�^�(�X��^X&v���074��x�v ��� g�?�fN���5[b5ƽѷ��1�����q�lU9�'iQ�:w�1�Ǜ	i�N̮�^Q� ������j��*�s�a��ۏ�(Z\�Bak�wʺ�[����}�E�����M��������c��ʛZ�/����>�,0�:�#��Es�1�Y�ȿ|\��n�	{���v��V���g�� ��T��&�au@	`�=C?����[t�|}�q_��kAH�ݩ�ZF�qd��p��������xyvӄ� �NOGG�c�e��@`�w��V�������y�>�����<�8&��ラ/�tZx�����%��:��>�{ 8ֹ���&Ϻ_#b$������$�YW�8� �y�1����i:֠t�۟��ɫ �<�i00q*�-���	���-���?�e�4��&����&��7�:N1t�8l=xM�hp�0Է�v��/��P���qWZ�@����X��Hj��-��!���G�`�=`"�^%�Fa�j�}�+��v��w��a���w�ڭ�5�L�x�-���.����̃��̯�0	���i9�7�P�(~C��]3^�P��=�!�I�E��$ϳ� �lh�J��td��/Yިۆ��/�C���ueO-xi��z������-��Y��W�=C�DsH�����u�ˍK��ga� Z��r���?s.�Ĺ8/�l�?����I��㠣��RQ�il������v3Κ^I�ϳ8��z��P8�H����
�)9�\��΀Q[{vn}��\PG>��d��BA�L���|���C��?M��mJ��[,��K����+��Rƶ���b�
2�`��cm�cr~̐�ݏ�����%��>�>��x��e�|�����kЍ��,M�}�\�����%3 H�y�[��jR���4Lfu���2}�{tɶaâ����R��/8�u���SnM�r\�����`"�Ǐ#%Vf[�O��a�7�>���h�d�$�B�t.�P��1��l�/����O�F�#2ݐF߾����D�׳,wc{�59�"�#�UȪ�Ԯ�uTG��Y!�^�+m�h�7��
G	����{�8��f��@N��!��m�Ii�$�U��l|�*(�=;�����k���,��ėzL��?i����u�O;�e�	&�A Pr���WMr���/ ���"Jy�| A�v[�.�ҧ*%�{TFL�ؕ�By&���(-N� -Nx�"r6{�{��f�Ǩ,�' `g��g�&�}Ё6ϯ�Qu)޳��dvo���( <jC�/_;��p�����:�a0����4����UOCcO�bf3�+��r���Ϣ���:��;�)\AR�4�����X|�����z�$��~�ch����!�<�8
�#��&4O����3�7�펿��bj�c����
�����0 �D׋T������_�̵GڵH��),4�$k�UDi1��ݕ1����\">qXJR��@ фp�� ��X/]z��`�J��.^i�S���G&cw5\L!�pg~���}���#kBI�M��_QM��ht��k6���쥢�)+q���w!g��;9�)Ku�Cu@��G ����r�]t�W�=��?�l�π�-�I`+^�4��J��y�KB�8!|v��E�.X��]�ܸ-�Bk��Z�f��
����%aW���r�[�h{��C��+H_;j��GG�ZUқ���VRqM���R�4Q�_ǐ��IX��K��<n$��^K��WQ��Lt���(}y8���,�"���=� ����p*wЮ�`$�8���\O���ʇ�~�8h}$�;?�?cR?��>�o�|���_CVh�QF���:�9p�d�1��8�s�ֿ�@bH�H\�-m����)�GH�X�e	zR���Q�����`y_���C4l�y�w���ACh�s�RIcv@�q^`x�#���x л������TJ{Mb\�NT{Nۮ�5��P��4K?�<�Y�>�>E#�+Q�xſ����^ߗ�o{��|��4�	DLJ2)�\ �A����1�̓ ��՚��Ne?�<����j���?x��p�i��~!D�!o�,YM�E�|c1�1-F���1��D�jk�F�j�*n0���'�`��3xeC#�Ղ�@�D~6�ό{~�ό1�ԩBSc��������S��T�ѓߤr��7Tr�yE�b����4�Ie��1��8�q
����ů��7�<�كn��O͘z�/�D�F#���N·�8;b"��}�bW���U6��82풥
��N�O�[S6��D?��m�V�8屙��	���2X:&_�Lz���������y�N����K:�*�!�)K[��CQ�_�&9
�1J��Eӕ��j����>�ש��o���R��l���V�����F�g���h���-+���>��&�1�<�R���`X�C��0����$Q�C�Ҭ�g-�RBn|���aj����q7a@D ��i�9��% �?��܆���07
����`��o<Ϟnn��=����=4��;Nc5�M���+C�H�?"�(n�;.1��~>�|�t����{pZ)�~5���5W�c��!�Ϊ��M|�]0���B��>G�U����3^�������e/j��F�4-�~I\�_ul����~�����_.�;�����'��{��������ج-w�E��J���&��{+9>���i����bn���پKD�ed*�ŸWϖ�&{<>���x �z���c^UL�
Sn�[��g���J1㤡|2k����<����)35}#���g
�00�n����c�v2��q~91��k�7��I��g~Td[̫4��Wu�\�/4�f;�o��ܰ>j�/]4�*�0
1_2�)�(	Da��9o6��ʋ	�g�Q��_v�=�y���e+0�Bڏ��}��[���y:[�M|1��+�NGUu+�����������=�k(�W�L@�l�FI&υ�!���Z~sB��֮�m��Etz/u�*"��ߛ�'Xc��}*(DѮ8����<��,�v�H�������Rt/W��X(������2j��<��D��?Bg��"��A���!s�|A����|�٦���S��%?�����;׏�����Eu��eSa;���� �!ii;�A\��]g��a�TF��m�O�����!�C��A��|s|?�q�� �8mr}zst|T�:���a>)�����:V���@L9*�]2˞��_`Wk�Qw0�(����R:N�i�Dwv�.��.9
e��wgo�X��2���+�ϳ�jZ�fU�k)Zz�l%�[�Ŝ�`)���{}�g����=Jmi)��S�JV<�8�?q�w�'�^+B L���+���B/�{���Umq)�K���(y*pn�"\$��+�a��awHa�R�࠱����K`dz�b�M�����|E�-M��#��&!c�jƥB!@k.�wu_2�<�;�vpM���-@�B��2�
h�����١�Y}�1��|��	ϓ�+�`˙lʐ�
%RWB��^Y�N�@^���$l��R
�<�3eZI�MO��S���]ԉx�����3mՕE3��|���̜��[�|�'.�NÞ]4VW��(�5��|�޺K�j���T�h�X����k]S@���и)�vu�Ӱ�l�-z[��{���x�[o��(�l|�����[b��I>5�yb���	�v�_|��I�9/p�;�G4׽{am�P���M�b@��X�,sP�Z2BUV�[�IǗ`&'�Wh�,k�r軦
���Q���ygo�-��<��/�'!m���*�͗Ѕ\%�j���_�$d2��4�=��4�\�"�=振$�=��G�F���۪���N���W����;�.�T������@�N���AܖJ-/��X��$�����2��t؛nm&1���Sp�̘�Ñ+.�ś���EE[YA+)���� ��S[��l˄|�AB5�G��NL��geꔗ1�ח [Z>x�~xB�4y�SU�4։�yAҮ�vE6m����Q�i9���i�K�J�7�?�]3�C3�p���re��J�R!�vDSU~AQ0��o Z����~���P��f��~�8�Z��!:/��G���� �C��R$��#����F���DB�'^uuY̬i��DN��z�G`�U�6�s[[0~P���$ח%#����,��ք��� B��RdWc#c5�ѳ�4Pۄǯ� P�ɚ�v�غ��.?m�I�;,��7�1��{lj��-�I���s �D�'F�����d�����g���1�^�4k�%�vjrB�<?��v~�O%f���S�-w��q��
a� ȈTR�>fΠ�dd1����ޙ��j2+���D�?�A!���[�+?]�L��(�r������4*�g�z�z|�eI�1�ۛ�ԛ�W)�O|����
I}�"x���εοM�΂����^��	?f�������f�x�b����]�6�~|�fRJ����[n>ˍׯ�V����d�9b�C��|�4�'����B3jaa!P�~_��!
?�5�4hLz��0�X�����:zy����sb��A(g��3ٗ1�W�fY��[Pb�������ӗ����Ջ�s�$H�7�����f�"��`ƭj��F/9��$�������.=�Aq'���X.5*G�����!�vƲ����"� :��Ʌ����VV�y/ϵ]����^:r�&�TQ�"I��F�H�4	��2�Dg>����`PHB���Ib�]@���aI9�5=W����8k�B�[���>˚�C�۷����Vߒ�fl���ٖ:coޖ��7�N����Zu�;�v��w?v��>�9��ZJ����98:��6od����������9n��[a뱤���弙&;����#v8��dK_������0 ��1��߿�Tk:�:���}��)�غ`#��A��|��;���&!&懏�-b�Lͼ�^v�����s�a�n2�8�R�k�[D�.�0ʆ��$Y���!VwȒ��%˭+�.�~0�� Y.���.���@����.]ɾchH&�,�oT��� � U`��2��K= �h�g�	��|:}�x��[�D���&<���RCכּsv���Wc`�F܁$� ��ˏ^~~�}���Pݠ?g�( �5��6#x�[�B'�c�2M	m}�����3P�ɭ3s�G���+��\���++����c'���eL95�����R�q�k��Ylh\rj4u_"zxx���>�p�321(9'�6�M3x0H���L%����M�:F|s<�q�'(���P�6e���;W����/�4�V��( ��R�� ��_;��֓L�Gx�I�I	��e5N�a�A 
�*���-g���tӶT���z?�'!D��Q������'���>˩�β�ư���WWxG��r i� <�遱��B�61�ɚ	��Ze�������{��8��Uw$~pISۺ�	�N	�z���N����h��z�ُY�7�ˍ\�ozXF��$G�J��kSE�E�������SW)��8fw	�d���c��a�Y��4�2�5�)�P^<D7Q�dC������Y�h�K�'���1l:��J�9�_��:kT�:�8�
5GAڒ�|�J������4kGU�,NLS"��.]K��i�A��)K��:�H��\��	N�i��������!�ׯ%j(�T��b�}k/�� A�Gw-!����ɥ؄��NCO�O�8 �*��Ű�s-`�����k�ğ�g��(V~ӵ�_#]�e�F��x����N�w���S��&\�F�W��4��}�A8���o�Ź��G5�����.01S�o2����>Sb?k-���1Ҙ�}1}����y���(�	�D��ɵ�a�F���C�9�i�j/� u0�ʧ��Cl���c~n��ˇ6�"��@Y�F�،�$����c��~-����th���2�� ������9���[
�I���^�N������C�ئ�_l���;��kkϨQ�]��I�QLu�G�l�I��s��YPI��Ԁ�X3{�`����Y�vh.� �ɕؑ,���ummn�N�6��l�.Fա�,9[���5�D+�fWaI*JmjEb�ymR'�@F���wE�k�B�v]R1;�g������6��7��2� �@zJޘ�Lw6��a�U4/�'��(ݰ�V�؄@��rHݾ;�t��A�`�J7J�����_�!sz�1�PXg}�r�LO~��c�~'�\,��t�S0�9-=�2Dq��nsX�r�~�������zm�H�DΊ���)�Õ���p��O0M����}KX�B������ni\�����TLg74pM���ثX�ƥՀ�^�r��X�����F;5L�G�WY5GR��uџ��������~w��#z)��\N���!�_�n���i�7_�8$�~ٱ6�,�-���y�俩�����y�	���������������%^�N���s^�T��g
q�l��*�*��4z��e"�.�H��!SWSf�D���y���R�n��Lq,_p�oZ����FB�oؔ�DA^r��ȯS�!�j(���q�Xq�j	�*c�g=�"mJ�^�k�ڇg�|H���? �"��r�V�D�'�}8=��^��v
����`*�jnL�|w~9^�g]K��j4\��!8�@�i�,� a�P.�!N��>���;��n�	x�7G���<��T�XE����]��'����A��-�r�j��~�Ӊ�O{�1삿8 g����}�h����/XD�p�Z��nGm9K\y�U�N�(��}�ڇAZϬA|E_&�>��n�EL�{A~�v��'/?�a��о������5X�&�JKlq��6�:e������o�S���MH�FMm��&�!(R��øM���3��֖��y[��� .R��0L}٭�ko)�Ȃ�r��H;��ypkk+�z�Y3�67E~���f�\jc2.�M�P�HU�PÛ��]��LџD��w�q֮> |�7�(So�Jf�5~�eũ�ڲ�F�N ڬ����%�b���_�gH��1�w�K?k�TUU)h9.A}��V���Ń_ɯ|�Au,B�Y���E.��R%�آ����,�-~��Q�Z�m�B�U����B'd7�/��ˇY����B���UەF2J���~ZL���_^^*麻��qvtv��f�^O������H6my�BCZX�����m��
6��Р�c�{��)�_ �w8���$���7��u�0��Q�it��g����j0t$��:���ş��y,�f��?2;A8��$0׎(ou|�� 3�)�˫�jN������	逍<�IҞ ��9�BMM}b��9R�Y��;�MR��h�E���?&P�RLug�*�
�ŋ"-S�-��5J��a�ݼ�3RM��x5J �_5��a�to
�ʩB*e��PK   '�8Z�ڟ.�M �R /   images/dcf4c277-9ca7-4718-9875-b39da06c9102.png<{cx$L�u��X�؍m;��N6�mmlsb�؍m۶�%���1�y���TթS��a�b�p�p   ��� ������7�O  � �J�:�ОJ}��+.34H��h������"Ƞ@�ب�u���*���i
���	��������8��Mkg����,�R��9�a��.�tX���<�2�����5a�{�$)S&P~Gw�&,)惤([s�̌bbb�������뷎<��;Nd�ﯘ�I�W9�oϭ���van1`6>��d BLyBf�ٛ�Ż,��ݥɟY<4�5������d h��VF�D�LL&5�Z�z*%��Gs�p���(`0��	#��uK���������|"�a�䅊\���^p�����#��]�/Y���}d��p� �!l|E?����X�;�:�fL'�6;���#h��K6�G3��H�~ً�ߦ��wSKS)�
�q��~�#�!|t���n���:��Ϙ
��?N{���'DX�D��x]�{K��t~q��!�L2	�񾹗��i+W�O���H2�Lι��H�1��v�6w�Q�-��W�h'�luX�P���^9_�i0Xp�W�g
 k|`W�i��������@m/���G�Yٛk!2�$}�菪��H"�G���?�V'������B_����BM��	�.���!�^S�ɍ��=�'�D��=��(����J��L���1���M���P�X5�H ��@S���%6�
D�ubp/���!�%��|������/ /3�A�0dg�+�m�#a��{L,�ɼ��f"����$�۠(�ٸ�d���p6���짿NP�����7 �(#D]|9��Ο��V�ǜ�������DD~T��֊���c����d�	C��!�@i,�9J'� b�ԏCQXFH�R��#��>�zX��+N�x�+�t�
����^\ cPȒ%�+�#�x��_PH(aFЁC���I�{g8_��4ɾ
�=�3��¾�$:Mމ�6�JB6y~����=�6�L�o�����Xw�r���x�����`�P�!Eȼ�aaa�~��e�ɿ4����ǋ}�7_��rv���?��6��KP����v&��Y<O|�G�!�<n���e�U�����Dh��h�RrU��B ������h6J+w!~� ��:���b6�[i6�qƼ����qǂ��~��Yn�"�U��`�:Z��}ۍg��,���9�8�I���Y,V�h�մ��M*���y�:����n*���f��	�&�v�zؖY９t�A�{�oq��Ӝ-���#��J�4�Mi,V����v��5�~�?1�/�Kȃ���Y�bC7M4-g�p"r�_�m��{	(�J�t��L��)�����ʴ��̳Ś���U�������Xõ������jI�:_����`�n�y�*�J�(��!�6������;)�	�v���|q�������}>���3T��ίW�tC!�M:�-��+�:]ӵ�+��i]0��`s�Y��?�x:C�QT��ȳ�'&���~T�l��9�K�| ?й�n�d�H.��CZP��!�L�B�I��t�����:=�xNYT����c$�3�.h������c�h�1_(a���I���Ϛ�x�\`������T�?�z��9��Op��0E��S���������)tZ��
���^��CAC��t'��L1����Z�� ����t����"�����2��M`>Np�Ʌ@P���аs�ֶ�_�g���e�����@_,3�Ҥ���ֿ�%����l{9�A
�����.Tj��<pB^�C?9;���KP�����]aE�8{��Zq�5I}k��+S]S�P�b�]}�� �� -����	ْ	��WO�*�.��M��;U��eM��_�W>��KYZ�Bz?9�E�[0���ks����Y��v�_���4�u�z+�Y��-칑�WU)�)�	�mFrߒ��E�.Ӻ+X��t��d&�(�d''/l1��Vh6��pە�K"Y���f�j�Z;_�r�}}+����� �X7h���2J��������o�d��Zhj�����Z�C=�ק�3Zao/t�p�}c�[l�0��b�M����u�����"���}E/ز�R���c}���zղ��L��e����<��0;�J��,�ɨZ��"�M�!�0����z�HD��b�qؐ�c�H"�@�,�JI��m�@�����\��$�hT�v6O���̀���*;/����vY_"� ޏ�@��Qd�A'W�#}SM*v▊	 ����u���@��Y���K�����wŋFy�|���H�2���W�ٳ�9�pQ��|7��c퐑�GQ��&}����ZE�=���[ 1�n���������NH4o �R�Jƌ�pP滲M�-�0_.�2��6��ם���h�9#��,�� pC]�J���s��z$c9��"�\�Cd�*�
�i��}�3b�*F�(�(���H0a/q �}��7$NX"b���$0��[�7���m�V��%0@�OɤZ���θ[��\���j0�Q$�{���wm�cM�I��'ׅ�o7�dm�g�`2G\��+<��ݯ$	?��/1�/�m�Ip~6.QRN��~/�<e�S����]�po��x�T�������I��Z�z�ӀkR40 �����o'i! �=%���<!
��:
R�Xoݥ!�V��`YA��|���PR9����d�5�
QD<ƨOc�O�"�3y��F�X4�χC~��N(��)�=`�uPf�V=_a�Pze��޽��4�s�Y��Xt���o���o�-D���Eh�J�[V�u�VB�3kk^��/M��&��ת��oT0�sJ"�W�`}7��|v�����	5i��P�}�O�D6Fe:Ӭ��LQ*�� **�HiA��D%�H�>8�b���D9�`���s�L$1(�,���h*6�O0
�ѾIР@����BM��;��i��M�)�L��gWi5��.Y��Ū����Ł��C#.��\�p2O��$g�������:�˒�m��c>�3؃���&WWW�
2X�G�a�|�I]�7U��:)�W#�Er�d^�8 �y�b�%�M����x~�P��f���C�0�(��T4�ᣥM�;	&����R�&(އy���Jiv��aev�I��g��nH�S�8���L���H�~B��")Ė���C�a+Yi`���+�sH9:�k�������LK�Ө�@��\�;f� ��e5I2&���`�Z޵N�������rz3��c�G6���I����/�I��������s�1[����n�l���o���
�h~$���ҹ���p"�E�V��}#�iO�����&K��W�����۶�۶jV������(�Wr�F����=1�(=!&�6#ب*�>�+��,�O�e�C�!��H�__A�S�j1�P��:L��!A���Ԣ!�H3��H5���p�[���)̹b�i?����	�{��t¿�|��y����{�䯴^됻>����&�팊��������.	J�=ׇa�Ro&��.}�P�W�pZ���L w����R޽{S�v�ׯ���cĵ�#E'$�&4d+���|���K4�]#�l���Ѝ�Qi�}}�j���z�끪ş��D	��Kz78\���6nT���U*����1��(�Wa�hT+fʌ^���,*�K%XL�� [2���56��{(���A���h���ſLS�H����Oմ$v��A�髑���Kl�|��/��V\���]�1�$�>�R���x*���-1�A������e�\���qUD�so��$_��{=�)_�r*S����ݏQ��K���EF�Bq��W�BX��ƥA,ƈc��D$~G�
�q9��2�=l�J�������s�|+�x��cw�f���\p}j�R�R���?�b��/_��|c�{�Y�@d�-���w_�J��ɰ�?&'|ЈG�8X-SC=����|�Q ����݃���<K��F��>��)CK#w��#r�5$$cQ�Q8�;=Aߘdl��p�T�H$Q��a $}��~����4<����=����.���L>tZ��tL�࠸�N?�=�
��Qr�T�v�=�[�����>�}��gs���r#`�r�[�էY�p�������[s����	V���L�6��^�b9C��-D‭������G)#���([�����C@�����ѳ�D�nZ���k@H�752�V�����r��d 	#��jyzv��س�Z&�	WX���1�e5��+�C�0�Q:�=Y�^��XL�ج�)G�����5Uo���e�[[�P�HrD֯M8�Cw8���4�[,�.�!����B��NCq��S�,�
��;�	��^Ǩ��)
F1D�{N�$u�1�9�~t|&c�S��Ь8�7hY��ĞJ���s�M x`>jj8��>s��%i�M+�45�i����v��������gl|���}�4|�lގƔCYYH/�0H�u��L�Ai���u�|��{
�8�`�R�m������uXݗ��������@�V�}aP��E�^�9��'k��F�;�T-�t,~�z�*26��XOIF��<[�>�C�B[g=�[LY?c���f��G@����v[�ۓ��5Ay��������,�Z�3���3mP5��_M�iQ��F�ʚ;*���&=l�����������t[h�L�����
5�2��0�����۟��D� ,�LkeXs���@�/G	��"�������0�S�c��b�J!I|�K��*�V���{�2�G�+�u��w�ĳf�����z>,�}}3rs��]��5�����C9�?-��7���x�c�~�	�r����tVi���؞��	]ϱ=G(�)-4y(�pM_/?R�����9���k��ؙ��t�����$ξބ��n�?��	�,M;�޾���A����T ��p�i��m����\�IǆJi�L�����d�����i<�Բ��XQ*����������tDMVŮ�~�y4|�z�oPB.:_�G�](�d�d⮴Fa�u�] �F$x���ʜ��x�Q�+�I}�U0�H�-V��=>H�n0&�2w���=�:�'���J7�{������ME��sς�H��o��ܘ��f��-������׀��̬Ue�Ƣ�X���<��hk�+)Di'�<	�����*��nv�h�I��N=�~k��/);50!Ɯ��: �p��5_�������3Ǔ�lp�&�5��!�;�}��N���l���G'e����2g�պ��ۘ��,͋��dV��9rR8h��L������Pm��Buy±����぀�^C�B	>"2<̄^����}�����H[�D�
B,�XAa4 n~��`��E6 ��$�P��G΅X/~����uf=\@�X��l���N��3J�b��Ad�(č��w�8S0�,!�Ѩ}�;Y��ΎƯ����p>Wk�q�'�O|_#����/qVumΉ�n�~�)EIz?:Nm�'��Qkqr�v�൯�Ҡ0\k�z)o����!О��(М܋`���(�p_��a�럈��tֱ��l�Cg��,�ק}���T�!
�����I��}�x3�~��/������UΕ���Q-F�~=�:S�X�����_�}�˩a���v/l���z���r&%5yV	.�Fl,n��qt�ޢ��x'�����}����p��_��"[{�	��Z�\���U����N�����J�Fǃ�m$��.�%�v��HJ|�;���ȕ�͒�Lk�H�϶���3:�G��ߑBJ:�"��b�}>����������L3�	�2���O�~~��J4iÿ�5|�MOw0�~�7,�^�>��:��ӣ풑uyS��v3��0UDO\�x<�J�p���P�ux.�2��*s�O��Q��b���]�ʹp},]'o�NKV5�B�kדB��ڧ"1 Vw+%�-T*N����[��`���o�;_�GJ*�xD���Ē��rWhF0Ƿ�U�^X�l���K��Wս���VwF!���������je�v�o���@E�XL�+~؄�Tu�W��(���w�������v���&�4�ˤ	��6�	�f���Lc<��']�	����~�d}8)�Ť�������j��?G����'�tDt���[{#c '�.�_ɴK�4dٴ=��x���l��J�lV�
uV~$&c�u�"'��ܷ�J]v:�p+����q5��rு�h��_�y~<��C�)�[�w�2uW]���'��x9Q�0�=��6���w7@��W�m����?����:�8AQ-�S-
*�?�	��m�o?0��'c������oͽ�6׀8,JSTcO �o�>ׅb���}|@c�
+4���*��k9��:ӏ�\8	��Df!d�����cs�}O����V'�0��2�]A�Rl�DŰmĳ��0�N̚���O�L��X�% 0�(,"�$�.)��I2�!>D6�-S��ȉq����Q�
2=R���0%��+H>���A�qL=�r��~��������54��;VNjOup_(��ʨ>���)Z�G����Y���v�?�bM��:��UY����|����.Jk�4��JM�P�����Sh|^8�]�&QT��A�,�9χ5�����3����H�Ј�Xс��������z�)lH���A�Q�W��[=�4�����a��t%��U���Q�5�����˽���a��.�}[���F�>{Gd����t$��{f�Uo#���j���h�2����nޥ����,(��U�i��%b�Rvė���I��Q�M��F^�̊X�1E�>�V�k]|ÌI�V�� ��9|��w-[���Wd��h8}�R<u4��>ζjE
3һ��1*띹v��*����$�Q�-"5�c��X�Z&��*���E�N+VY|?�QF��F�ͣ���[��N�0�KFx��
ai�3��0+SB�?jYKj0W,��z̯�AY1F�,yh�Ic~R ͟��G�LջC�y_�"*�k�y��/��A:����Pf���(� ����.��4v�E㷰��Y9��XS_�
�?����u�ݿF�ia�"�:Mgɥ�V�����pn~Mo�܏G��!i��G��BI��L{���
��85Y�������ݘ�xW�O�$�"`��R��5����+�v�uc���I\�ټ#2=8>"�|�iCp���T���(+��_��@'Sw�X� V��|z�f�ҋ>۬`�.�?��w��pP�U��B� �{��ƧO�ei�åYdf`�#]�}K"���l�
A�5(i6�|$���ъ�r�qHq�~ƤB/2,썖w���^<{o8I��zm��K�2��K'���1�5�N�+Z��s`�Y���K	�S��	_�i�p���ޝ��w��#�ԋ!2$���cj�U�o��9�Y�RY��pϗ���ܺ��K�Q"�vc���P0P��cI$˸�ۓ�)m4��ݽ�|�j��/W���3S��7~h ].�|�8��>�vF�)�;;{s�h�)��9�1Y;�@�t{�״���Jl�si�h.C�*7�؆35Ud�y|i�y �i�2+a�&%�VՔ����9:.cZJ��p�=��a����鑿Yj/"�;��f�P]�ys-'gZK�G�����R��X����r�X��|��U�]�$�1ُb��\�
��d�j��㳚��5>g�(T,�9��@���Y);���I"H����°�Ⱥ 0M���-d|����4R��*R�Zvte�r�sێ����0%�_��6��1��Ӂ��2��\֫�f��I}lCh_EeT�%`2��b?2O�
7�EĤC�w4YWt��iha[m���N)"y���!i�CH�N~ui4<��}���WavV�6��֚�Y}�ФR&�+vG��W�jNF��6��iH^Q�$j�`}���d��L��
�hV���a_S]�zf��z�/�7�o���5)��ྠw?r�Η�]d�¿58�hG��;�GS�3QI�1���*&T����l�H'�+3-��w@rq�ܳ�F�F+;74B��c
������l�'�����l@���_�����Ç��P`�����9���D����*����Bf�{�	TSي�1h�9$���k��	�t9�S�9ۭ�� @�x��Q-�x��}�ʶ���J�����Z�9h����*Z �=�L�K|±/�jI��+IAmE<��c��2���<��?������ʦ�p������z�9B��=��֭04�P�S$�&X$W�J�^�WWBv�n^���M��&٨��X�,n&'�*��]zS�ɟ��%�e�6���.���Y�v
Ң-�(C䉛���yk�%X�:_�/O''#���
�A���੖\}c-�f�EH��%B��tr���c6��ˈ�����*��� �ZG�'>O}��nج�(x/������dDiGZjA���5M<��gh�\�/�����C�����?�(��I(��bb���ZYNDp�9UQK�H���e�Yw7�� +���3��	��B)CF�*�VZ�H&�)��nG�b����	�����=%
d?H2��N� ���T���(�ƺ�p��+��;�����b��
�<���*�Ķ;�P��γ�bY�N�������Ŏ?���7��瞧pk2��&-$馋]>~�?ut�8�E�`*+0���;_�t-[>=U�֐�ṾC�+�J�X��Ղ��Q��Z�?���N� ;"�%���%̒�*d� zc�6�3e����L�LN'�c���!7J���iN��QR���/s��3g=�yl|�i����&�)���V�r����N��糦K� 
����UZx�rU-��X3f��Xo����J�X���e�v2��������c�j�3������uwH�`���p�EI	�پ�A�n9�Hn�#bi|���]w��;�qy�b��A�&�@Gu�����I��6��O����a!R�&;2Z�9���c�2ߧ��T��������4?OaB��V�z���]�1�|�_���p���	\�j�ۊAC�_n�x�-��A�~D5hA��1�y���)�|�*8sT*��[+I��9ϓ� A�@�����JW�@e��<&�i��K���p8l%��Qfe�=o�tD1�7�ca2�fjiX�M͂��m���-R���,^�&�k�s:�jJ���?�8��e��_c�������Gp��F��н8J��~���U�F鳭�!kn�A�i!��=�a-��<��R���B~uoϑ��N�e�I%�k��\�t���A��Z9�2�:�Y��B�c/�0v��z���`������ui	�ΜN�'�
-�ذ��P��O���b�K�CW���"��2���:�G�E�?u�N��+���.�7v�����n�f�+����*� %[n�Rh%�󱃯	������r����"(8�.��~י� �~��ş����13Q2m��"�߾��Z���Jh�s�B��(�.@+�=�cuJ�D;�nw����h<!�"�!������{��x~w$����z�^;�D�9�����$�VC�5�R��bk^�_�?��0��8��9ǃk`�����i�W��>���U*~Z
j�sd��h��a뾽�hB?E1�d�	ؘ y̌��F��@��B�u��H,��,�o(�+�fH��#��dR�IX���=��.tL��&�*�M6]T���1��c��1��\���,��,�ϔBu:��Y��ֻd;sp�M0�Juˣyx���>1O.��@��b�}q�(8S�w��Z7�/pw���+>���l�'��\^�����M�D�F�C��k�Xw	u`i6~\YC�NЫ.�@D���r����@���p�2&��BX���Btƥ�S�� ���bTZv�~�'�٪���{�z���}<��_�h��#�n}-m�y�Z� /Z��L �h�c0ۓD}K�J�s:_��xy�%���ĤhGx����h}��\���<徉�u����W�J�F��BW�dX獣Ӛ��`τ����UG�ùNf��a�;�bks�3�J�N��Ou���46�z>w�˞aW��Lq�S���W��	!�N:������k��4�����{��:�s<���Y��E �E8����8�F�G1uLdpT�1ʊ�N��Rk�w\�>�Z\�hu�4	�gQ������$ɲ�(�1���X}�/�5��m#c��R�9��-2R�E�`�1�ҍF 'l����������O��4��)�Q��Te�P���פ#���<V��U���k��X�Ns�%���t�P�����[�$�ʓcK75j���J<i��)�w���A3=��;eu�HИ�x�{�-f��=E4�J����~�Z=�+���~q�1�Z���D�ۍ�y����Uo�f�t����,xxxAϓ6��p*cmdR�+�˭�g�:S�	���r��M�*�#��ɉX����g�&n''	���d
�1DX�#جo��L�F���O�YS��⦭c @%�ڟ�.{�l�^$��R������vuw���.^yITF��3�C��Gw�ꤖH0�B�nI���@���$hh��:�4{5S[59,��;��wNxXvÌ~�����?��q_����z︻�ȭ������~t�	�h�7���[�����j;�wP�*'Q)^��W��T3%����둭/��ơxc�Aͼ>؇�=Nͷ�Tθ�m�7�V�\�E�4���x��W|8�K��n�?a����~F�Ap�����e��R�E;ERÂ��V)υLg�B�߫��m���Xܝ��@$;�����m����솋/�&ml�k3μ�*
,LjُK�`��M&Q��/�W�Y�lZC[�? P dXo��Pp��<��:��)�Y���t:�)�&�� *ؒ�����i��{�c��:�>5�i�&��|�00�Ϧ���(G�q�l��0߈��7չb=7CQ��A�E�9R��a�lr'����xQ���`�~�\T�ËE���J�r�ڒ!�2��_�ƫ͹O�d���P|�R�Ŧ}q�m�T�6�޲��Ao7IK�{��ӧ��yk�|�5�n746/�͔u-0���`�[�Nd�dƃ)�p��H���h�(�Q��w�Ӷd�"���8f �[��g�PDͯ�x4��`����m�U(W:�X�(�(��>>w�]��'S�z�}�*�	cl�:Ϭ/(8����{,�Hݲ@�6��Z����F�����VȖ�aT���s�/�+��{LI�MQ� �Xw����K������s$���U�2o-�Y��A� ���JQ٘�z������ ��
��O����ӹ[H8���rժ����E�P�I �<gP�i�o�"+z��zu��V,��i ��8v�����}�N*S�=Vo�	8d�|�W������}t��:�)�}�P*��2s̈́^c���Y��9dU�O��V�Z�L�
������[����xq����[qr���ɏR�r�h�>�A	6�
�=�z�Rp����2�̡�
���+S��o�ޕu�{���V���̈����N�����������r��+��K�n��T+D�%Zu\u�A�^^^/��Ē��%�<�^ʿ��r;�-B�^/Zm�V�(7=\ցJ�����G��w���=E<NK%>��9��mՔ�QJ�촆,�u�y���a���=������$B*~L�	i#[Y�(�=9�J5ʆ�F���E��1���h�x�[2��%�?�����Y����ܲ-�'L����8�2��	mn��$��;D�Q��95ZQ�G���|�5!M���w��v	�3P���ߨTT&P��yٔ�ax?��#��%�[ݮ��DU�jiO�~�Kf(+|�q���A֧k<yĝ�nw �e*tI�z�-������"��w/�s�Ou�8��u��O��a��䜰�j�o4+������1����_���H6 �v��:=x	�;g�A&�C���CW�h*u��?��l̼ҫտ�a��=!���	�W/�r�9���_���/�	v)�������n�0��|�vcq�s㉣�݃
��P�{!I��je���Mʹ��knH�Y�0�J���a᲌>���d�,�V|�s��y<�s��M��RP��9o�+��1těW(O~�P�+�0���!3]AA�o����H�F����Yu������eK�]����Ph"hT͝"�V�j��>q�߭�8\z���w��q���^��w��-�?�p�wD\o4��[��/P�f�nd�/3�J��z���4Wk�T z٥0��jq����6J�Ū�Z<E�g�X�'L��)� ���͗�J_&-Ǚ)$����N�E��b��� �S��#����{���|�n(ήDa�IR�N�"!m�M��V,@���t":�Aϲ�y!��؍�|f:��e:�4V��:�7���p4s`g�沀���D]���o-�6[��Z�<>ޔ�ɣN�й�@�y�5�]#檦��CV06_��w���)��	�8)���BCW�t�5��%�n
���ٙ�{�]��~
���[���
.���۩�q�E�@�a��.S!A���Tl�*�9�A�7i��E؈ �:O%{���tE'�zc���������5eGf���cP�cS�Ft�|��I����j�w�\���M����k�T�f�����/�J �Fv���<��p�nBv�<6�����]�_� ���Ɛ��i�c�K^Q ����@r�:91
�0!�3Y<b�2��7���Zn�xt�N�����~�:��[�Z�d� �p�t�C����)+��ZR%�E���pgwO�fȗ�B�W��*1��5�Vt��F�yq�Acp>{<����@X�h ��>ydeK��M�ޮ������=�L�y�W��n�����u}�D���tRQ�2�:[
����T�'�
'�c�B0���p�)��S,H�]>��Ko�l<>��r�	�9��P�5�8u��j�����UZ��C�1�KZ��<$$7Qr���|͜���?��`��;~~T�΅�]�26Gy�i�t��K�*C�M�[J�'����3�/���2A��
yw(G��N�Arn�KkX~8�i�\7�윃iie'�u���-|�=�����$�h�@�(�VP~���$��d8����飰)�g@N,��"��� -��`�r�c�����a:�W`�? ��j� 0�)��l4��(p~��o���bs�61�Վ���_�и: 4_��@�`F`��X{S��	gOǌC+����W��g�����Җ���n��N��Y?��������3�=0N��;㱈��bLY�����F�w (��9`���,����f�w�DpD7�fJ�A�>��I%���d�I~,�'u�� eEH�>S�]���U�$��$���3�t<[g����ޭ����'���L�y�J�FV�s��#:DP�U``�3����#�V&��G�g�u~V�����[��EF1�(9M1{ߠ6*���Y��\ѻ�DƯM
�}� [<����æ^���|��8���h^�~I�E�|�,D�K������9`t��I�l/��*�|�7���A*c �s�F�}��4�qH3	A�W���Z侐�c��w#�I@�b �p�xc"��I�<���N�z'[��5�(4֞����Vz'f����m!k�c��O��*_��jz{�]w��]��C�����������E[s-�x��P*���֭z*�hHȠ����K>ģ���]m�Ay	~�(9�᱒|*�78w'�@�"�=x�c�{���Ud	w��Ѫ~�^�FK��/�������?�m8=⶧vD��E�j��8u�>Ʈ�Z#�/��n����$���'(2a�/pF!�RM���a���"�T
Y��Go%�?��0�(���/J8��{�P�xHzw�QF�	yK�=vrd �f�䟞Q1�����z�]>yb�D�H(`��T<bQ^���6���ses�q�������v�"p�:b|<V-U����x�~z��-�8/6~(.BJ��L����lpVo밽���3���?-*�9~�PSɆ���.%v���y;h�7K�ɫ���Qv�Ӥz��P�$�ow\�Ni2��<ݝ`vJ��Qs���ó��,�;&$q��,1QdF�i�ZQ��	����C��E��ͼ��z�Xb��F)f�gb�a�ߧ��j��H�����PM*[����*�L��?v�fZJ��盽��� T��K��?o����b��k�0�$P�%�������=U��ͬx�\1F��>g��r�r�pĠ@_ ��z�9�㯹�A���8�e80h{a�0��̟-��,!�ifؚq?4J�Uiӱ鶔�T�=U�I�LdjC5��'�uMS��}+��Q�G.�_d\�"�k�
���B^_G�4�Sg_J~���J�B��ggY�u���l*��sjB!N�E�ʞYD^�jJ`{��;� ��2���������m�v��/H����jWO�dW:��z�>|�Q'�Î��_�k�~�a�L3윿��ݘ%�gr�ueӘ�d��*3Z?I���d������4��	��Ĝ�Z�eX|vv6���<�{���&�6JHTR<�@�&�3�v��Y̎�#�
^����J�ԩ���.	�8��X=ٍ��4�BS�l��_T]��x�$&��p�����6�1�!�x�B*��L+��§��Ժc���p�g����+��F����.6���T����؎kۗ���ֹ�j&@�L��F�߃�2�]
S�2��(�1�)��ON'Z5��^�iM�8O�� 33cFh��Ŷ=om��fR�3�����nT�t:ݗ0@@/�h Ne�bY<x	�JP��jܼ5������[��C��V�-v�M���h∐�s�I��?.|�8kS�8��6�Gxӻ,�_�q�o3vB����z���#����g���N����_�+u��������(e�p���r��ڝ�
M.�Ѐ�7����u�ﳧXna��63�3;����?~w��.����-t<��S��HrE#��(��]����y�Z�Z�-y�BѐIt���+m����ԐE
�����$�Z�3�,\�_��KAU֚$:^F���b ���ْl�e�˴o��C��@@M��GnߞT�3��2�QV�"����ŻntT��wW	�)`sUҢ�u���e"����(�ŵ�n����6�����"$�r��n��--ǹ�����>�!��p��]�mu-:�~9��V�L*�;אq�G�Ϟ<h��|�m���������wض�=dy��_�kMr���uej޽.;�:� X�f�s�#�����E�,�$P-[�J�f ��n�NӋ�z�}*~(*���~��]���ؑ�)�Ð`�$ �����x�laK�s&E�֔Ȭ���t^缥�s��,�e�{OI$ͧD"d��,Ż�����D�c<4���ݝ��Q��{�n�:Y�F/X�$Ҫ��$G�x��)�iz�P��K[~뽨�z/cDP�ء�p����﹫3��$�+ _�>��3�,I�୓�\�8گ�(�~�%B��j����TA�@����5E�)*�	��Q����*^��u�x}6��_n����7�XT it[q�ˇ��}�\��1kl����@�`�O�\l~d��8�9k8��y�"g��3?^<$0��!������q|�z]6�\�D�
㓕��V�ݭ�c���O������I�Z��+	��1��8Ϻ�bdJw�7F,���7|.�{:����@�B���E�	�d�RIz���N�ձ�4�3�;���it$����S�|Vd2�S:}�P�bG�"?���]��I*G�^Dc�
�n��u��L�\�&�5Z�4����� �����j�s�±�8���ӿ��=���_^$��u��-� ��J����� B��R��Z�{��	PDi�@C��	�R�����E[�NenƦkN$@��}����B�\m�K��y%�َ�W���=����it������LZ��`q�X��y�w�#��ƾ7\Ge�U��C�bM��.��\oqf�s�H���C�铎��щj��g*,T^�M��*��~��Z�;�˵;UP\�!es�^�NO�[�c|i�c5m�� ����W6,��i�Ps���/��!��>[�i�&鋹r���)�+m�Hw"�� K$zk���+�p2\�?�sOGl�a�B%H�oZ�pK������9_�����/�J�02��X~sb�%&�^�9�7���-*��ۃ
g>+���g LG_�{�������O-�\	�-���];��W/~%�4�v����q4cZt��^�|��:yn`l��4LK[(�� �@p�-�#��do�i�ȩ�Nv.�7PG��T ���R�z�����_}=�)��k���e
�����LaeN��f����;YZ���Ν;����_�^�~�qXX�y��(X�����L�:d#��tr60�����h�6�,�D�R�V#e ��ಖt��V��J�x��)F��lS
.��3�M��N������}�����N��N>�Ak��ݚҿm����%K���4��Ν;�QS�^�z!���'O�m�����W�~���Lc8Sr�f���d����/
./����IHHp&:�^���Iͅ�c�x�E��K>�w�������h�H�;y{�v��d�{~N3��+i_M�.��Dk4R�=����hO�{�)}.��ʨ���II�4��R�Ւ����j�I_�@�'�~�ihϞ=w�Y��? >���W�[�f��p)�l@X����Y?q��l)>$��Y��nA�跗����m۵,<f�~;XZ�����k׮��\��suuepGF�!���7xJtt4KLL�F�s��B�#�����1ҩ�󌋋�5㟿������ￅ��*U�y{{mq,X�]�r�EDD��t� �_���FHX�D_{��u`�I #x!b�8�nt�S���B���c...�������s�P��"E�\;v�����{�"@|(�'����S?ٻn�5�Lɀ��k�'����KS���ٳ�<ݼqW~�� ����� c͖��(��K�����)9r$�O?���N�u���̫hѢ�E���?f%J�~� 0:A�K�.�ӧO��7o
}8C ���3�f��������7�A�{��{���=<<X���I�͛7�g`���̟K�h��3N3��w�` 9N~p �0�ށk�ʕY�F��=7x^�V��޽{��Sv��Iv��� �uM�4Y0w����~��F��x���[�Tt � ��Y�ʕ�R���ѣGF=<�Kg�Ҥ���nƸ8E�9*z0ep_���S�����K񓡗�9r$�����0����'F!��ݻw�ك�����!m@��'�N7˺c�`d`xU�T$R+	ʔ)#0��ϟ�G0>���K�\�ƥ	�7�p�ȲEe�� OX��"I�$Ђ�h��o�e����3HZ������� ]b�s�α�K�
�ą�ʗ/�a���_d��mJ�Ȕ�����Ŕ���+���ƙ9(�Ξ=�b���ݿ8��y��;��I#�b(�:���n����d�s���#���*1�J��թSG 02�.��#.];�x&�<��؅��8�-�a��9c�W�b�`b�W�lYP�鹱�� t\
 x��	��I����$�
����KY�J���{����Cu��f$u
�$MJ�#�=�Y�p�
��g�+�@G�b���(ṁ
�BR�-X�|��중�I���+(�Ѿ7a�-(Q�Pp�h60/��ÇtJiz�խ��P\��+ �jf�5{��+���k���r�4h��N�]p�8|����I?��:g�v��e.m��s5ɜ9s��Çf�1�P \�d������ց��.]��!���Y��p��ҭ[��r�<M�j�krI�����/9-�@�!����! �J۶m9�t `��
f��ki}fG�[��s���Y�0a����x�?a���;t�p.�� ���)�ǷZ�+
��
��0=�A�gʕ��q�o�R���z�ܢ��ܨ��Ťg�������]�<�T�v�d��²e�/^�:~�+Vd`�\U�;?�я�)1��5��3���v)b J0~���1cư�W�
L�Gv 7�r��7�����!���P�}��G���ۂ]��P@��/^��TdX'փq���7�r�qF��3W���ov�&�"�H
xV8�-�6m�~�ᇷishM���g�Ӛ��3����(�oFsA�W(x~ Q2�=}�T�����H%x6�k�? ����c��UjT*7�
K��;|�ȡ�5��u֬Y�SqK��ւ$��t�Cv���b*Юs��cƬO�L�^͛7���_�B/<�|V�X1���'�Q����l2�>�T��}N����]���$1�/��&�l�	 $;.~/�l����F bN����?���'�b)�h���&��ao�A59 %�06�����������=��Z
�w���/���g�3��TA ���=SC������] D۪��̢�+$���ٳg�ĉ9 EN�>�:y7�{F���Եq����&�I-��ޖ���z���+>�ZJC�*r$q(� �9�D͑?~�ٱ�o-6�ʕ+w�N|��@�"<x��:a=���ܛ��GF��,'Ch����8f̘�8��X��^:\eF�F� �d����7�8Nİ#�C	�[+�P+��j�J�Cp@�: ��$��ū���`t��Ž����3ą�����������S��������/�7�|#�!�D��/!u�x�3D�4i:�ԡ��B{T���;�� �7�`� I�_"@d9�S���'�#ǌ5Z������f�% 6��7_��������\�5k܎-]EGV��D~�V{��(��f`?���KL�:�gz�$��L ���+bp�ɵ��-�!����!"�JP���G�Bw`�X�m�$����^r)�{^��a�p�ũ���)��QP����V�* �0��D{��y��s��UP\�p�{]A�ޥKa,̅���2<�`1`� ��<wһ�l�5�  �p5�uq�t�Z�&�5��2)�&s���T��� �K�'�h���>���*ea�;v�2c�S�1��xV�\j<.����=׃�`ߑ�� 4��*�h�����|]��t�BmrK=�:�k֬y疚���ڠ1�x[nq���J�$S��O�`�%+x�d��9��hp_�
���y��$�`#@/^\�THh���:L�6M�"`���Q�V-!.�']04���c3g�dAAA a ���+b&`��D����я���o������;� O/�6�.��1黪$����|D���v%�Q �?8	`lR����S��X��L���)�cŊ���^}FnE�)R)�"ϟ?�b,Å����^��]E �`d����=�4����?�r��I�Ӕ�A0�5j�)S����Ǣ�y �!M�1�j	1��f_�����Ѽ  `6d;Ͽ��+�X�L� �լYSp���`�G����k0D�ḽt(�ɓ�\ &�}ǎ ������y;��>7n��`���������^��a�����.�{L��H�h����$�D�n�/�Q�j�ڷl�T"-��m�Y��}��Z�'�"Uj5����E!@�}��[��|��c9<G��Di�;�<k~�r�,�f��Nŭ)@n7�Z˖-�/.n�$��1։i!���)���y��}ɒ%�$�l����B�?1ꂭ:n�A`W@<N�8��_�@��� ���޽{�Ǆj�(N��1�� i *"Rٱ
*�E�1��$е[�nBD����?���={�`Ё���%���*3 lW����TH:W�v���<7�=�BN cq��)Z��X�\�vM��4��4lĄ�C'��_�&[塱��t�"�����۠���e�LM?HF)����i�;����4=�9�nY1�y��]�j��`q�ŉ-y1���0�J˽Ip��R�q}2
<\v���N����ږ����  �m�@�B�`�gP7�}�"� (<��a�3Bo߾���㏂����?g��������
lPUQN!�t�0H0��=$
n�E46�� �ѣG�e*ś�%g{{ OI���S ��D��d�	H��H�7����  (��$W��YJ�Q+-㥷�(A��r���/{�r�����:ʧDFj)��<O���������4��5%�#	�Z��
ߕ��:���:��'��60�֭[�~���s���A��i�~�I�\����	���Ǐ���봌��-$�@ ���
��Z�� O"�9�wc���S/N�����Ў�3J\(La[�[�� 	$� �4�6@�_~bI ���L�̏{<aސ8���F��{7R��70׷o_a��������[R<��w�ɛi=+�0.��1b�`#"��%U�����~:w�����b��n@ȕ��CBN~��:v�V�� 9f�1#��U��t�_?����~{�+��;lڴ)�
^;$Q�q0��@�;d�-��9�;O��&W��!�Bfdu�A\��S?N� 40θ��	�|5ڂ�c�8��?@1h����&�i��	'|���6B{���B #���4�	�$4A��s;	r:�B�م�2 c���i!w���4N��$*�&�<'���b�N� �$���mA�/���m� �~!D'Q�d+Asr�&M��y�&���� (���y��4�޷.�`;!��5���L�V��j�X���)�N�dZe�܉�u�J��qz�y���?���;h�U��<)��(:����R 	0O�0�@��1#���Ps���`�P���<P�8�C]�PHHȻS.2�b �H�$��y��  r`� 
�腋'�Ԁ�_0z���o_�K��4����8��^K0ރ��vd�<Yޗӟ��Bu5���`_�.�H��	�L#{�hЇ�8�~�ի���O�	���2VFۈ*��R0���ֹ������T�ps�J1�x�b�m���Y�\�֭+���%�k���%��S�ڍ��21�$((,�Sʳ�[�l���`��&!O�M?�G������)���ߏ�8��y�����ɓ'�Kؖ�\C���`�pS�� �d�燊	� )�Aõn�`�`�|�`��I���$ �u`CR�`���+�pH+�y�Č���DKAg	^Lmڴ<���
�aq*�}x��Z0R�s 	�Mk׮��瑫yL�r�J�Π)�h�v��$�B���3���zr�p۶m�sCRp�	2R7� �TN��JxCo����(E2IRoT����5kV�u��םE�z��e�jrq��+�'�v�̑��<�� �PC��Cғw���_��/NnH��9O����S]K����Σ��ψ��$ ����|ذa�k)#��M�\y���2`<0(0d��r��R�*#|(��b��:X<�3g�<557&s;TL�ƍ�m�C�I�	��xj�B|��������yV[�*p��a!s.��9�H� 8y�n�+�^��B������jI��מ�sф<�:S�� g�~���RDҞ'�h����־"@�J�,jW�f�&��icI~��!dW�]+`���[ ���I}�mܽ�K�#�%#39:Q&C��gUY4�<1,1�������v0Bds�i$��?xI J5�N�w�9 OD>b:�lZ�]C���#�/_�,D!s�Ť�e�hˣ�q̙��al�)�P-A��d�tٸ����������\��~!��s��R�}`�恊cC2�;,��N� "���IOH��%0X� ֯��b�āk�g��QX7�� 8����Һ"轑��9��� Յ��z�� �7pCM ������I�b������"@�H��jV3����l%c�^�\L�bf�7s��)������2�5>��P��̨��V;Gv9{F,���"=yW
\��s��A��*|��I?`^(��3.^;��]�*|P@���`����30e��rP� �y�C���I ��ŉ��y%W�T�v���1WD`t�rƩc�s$�]���yW~����^��+(Cr@55�r�@Ui��/��ā�g�Ś�Ό�JX3�?�kR��w�a�&\���L�^K8T ԓIt��s�a�Ff̯z��T���d"1��J#�w��MM�4n����֥�!�;��i�1�D�x����ŗgϾu�tQ��I�I�X�3�r�	��o>7���`p�x���ƜQ�Dn dq�= ��� ]�M���4�d���ڇ'���!1���Bm�{p|ƙ��p�w������e��`p�X�Z�w^I�h��h�x�qru	�k׮�;�L��`4�����J�fK:��ҟ�s���G`����4Ǟs���<����ā{	�t��@;���Ŕ�M�I}kՉJ���
�ҡr��ul۾��QÖ�o[۵>���i=䨒�J�^yx����1��\6��� q^��J�!�3��DuRK��2N���Cpu�h�#Ɖ�_0T0����m�z�7gܸ/�������)�v�FlxeF:m���LH���;�	h��)�:1WH��O�p��{(w��m�>�$�;�a?;ҕ�u��G�"R���RXs�@D�������/H���0B�=GD�Ċ*���~&���[�rH]�*��@Jfkުy�I)�t�ٶ�N��W�$F �>�h�E�^�o_�%J3a��zH('(������ # P�9�����I�]|�c ���	�>�����1��1y&S[�ʙ;?�s��#�:�K�<���1 )�� �$��̉���mŖ9��6� �{{al��PoqK�ԓ��2`�ํ@ˤ,���Y�O��{v�Ú�#�P@�v��U�6l`�z�}���It%�v�옿�A��X;� �-!�ʆҏM�����:�>h�{s��U�q����VOŅ{-�2�U>=�j���x99��� ��7Zs#$"T:TBp�ďL� d2%#� )�/������3͔��N�ܽ��	0@.���G�p��
�)Rj <����2�i�/��̊���Cj��{@ ����:\m�kw'���sz$͌�!+�r�Zcm�>�w�}xv�ܵ�^�!y�o�	�y&Id�I2�����c� �TN�~���,�7U�`F2P�H�4�W��ɠ��}�VԪ����PD��H?.�s�<8��67����^N��=�����iCr	����$0)#6�Ŝ��G�����Qs�Gn�@;�#-D�/�� (���u�_����`Ccx`��n�_����m��|�K��yH���} �� ��`�u�y��*�N22����cI�G�s�3~�ʄۂ�9�O���Aߤg�*�uլ���;Ȏ�����������d6��H-S��]�U��ݷ�$3C��
v?[_؅��T,�R$1���D��P|e>���	&�L߹�_�;w��� 2�x�?��{O~眽����k{āfA]��|I�.]��y\�.}���B1!�i{Z�8O9~ڿF��11�{?e0�/�C$
�!k����i�hV����3MA�]���ВJ<0���a���Ec���M$��q6�E[ܧ��V4���g�����LCL<�]qvR�M��o�P���o^�����W���9)��q�$�.t���R�J�@�P�n<�#��� Qc\�1��>�����!.�&丄���y�-����r=����.j�i��Eef�����������}��e�_\����_`���z%���V:� �Ph������i����g�K��Sqy�uq�IO���!�hHJy�"��4L�Y���9��T;ĵ�    IDAT��<B��!&JI(�j=����-�YEο���y�Ӈy<�zV�?�G�}�4Ԧ�s_��[pL�V���q���$�Q��|�)����3=n���>4-��IÆaBvB���uֲ�M�͊"?���t9�_�΍/��vW���,�(4��,!�2:���j4<@���%{o�.*oh�0�y�g���1mr$µ0��$����4j6�1o��MEn���L�s��i5��w�i��vGRk��`B�%�^�0y�����5���*r�U�-����3�1U������\�;�����{���U}�	�����1P��u���S�;�\n9��c'O7�]m�?���#�}T���Q<8�[}y�Y���CVe�PIM��B06�A��1�|�������~��2h�d�x�z�v����Q�CCܯz)�%p4ʉ�h3��	�����mx��ޤ��ϙ۳ւ��ch�{��@h�ϑa2�)�����q.���S�w�\��+��j����}�uk� �����t`V�+'s� �8�*�Y��� �c�ws�E�������Nmּ�|踔��j�M���=w�ڵ=��im:v���
�X�z ��J��i_�޽{��V������x��5��OC.:��P�V=k�Z�qu֩�y�i��(ǰ'צ���ylJSS;����	�J����{�=3[�pQ���מ�ßY�*�1>�:7M�s|�Tɕ�Rj��xg��Ȓ��g�yo�M �ގ\%n�c˖9�X�ܨ�uDޞؓ]��N޺���!G�A�6��{���:���x��,�/n�N���o.!t���k&����vy,z$|�����phl:��Xbl�����ACg��I�;|o�[�ә>�_�V�]y�%���Ǣ���͢C�)Q�U�
�ʷT���A��=�N�|��sN�e��x"�*��T_����	��ۑ���nΞ
1�sB�Ȅ��ܓ]m�/G�F�/% ����d��:����yi���d7L,_P������ȸ*I����
J���o� ?S/Ǟ>�ϵB��gAU�w����O4*�.\���s���R���:�O�IWc��<�^cEϻ4�dߟz<=FE��x����nv/�2�� ���B��9�n� �=�*\o۶�A���S�x�i�����P��[/(*,�����-Z��;bO��X���n���|19�e�e{�*8g�4�4.��^�ގ!��G���t�����IMͨҘ����ַ�D]uo�mO�ә/�K��C�NU��8V�����Z(H�\It���i����y;��Pʞ���cOR�"A�[>\�H�8��\B*���^z)AR���ޗ���λ#��;�}�Q���ɵ�m�roQ$���V5l��=�&�ήG  �2Sh4XG@W��sK��t�Uu�a���(t��F��A�ؐG�_��$x����Dbh�}Hb2sI��i�h�5S�*�VJ�ج"W�F+�9VJ�+��k`��i=[{�?dWUt|�\��zk�wU����m(=/�u�(����뢋.2�˸�?>��sբ��� vw��{��]���5C��.;���doY�pq(���r�hФE�t������C ���3fL⌜"wTp��_T6ڡ���}6Z���> =�c�3��z�iP"W�-h{P :��Ms�>�����U	=wd��?�p�z�(�xMc�v��t�_�+�}�5( �ִ���Y=�	4�Jڲj�pǎ�/&����zw��2�O De�b��a��n.W�:�$1CxOv���T$��8��E��{���'��+���yw��&�0Q��MZ�������2'0���.�m����x�Ep�H ����a��Qca�Ac�4��]h��=����Y��<&=�*5��#X���ABύ��{^�Μ5���O�r
2ꉔ�Ya����&��>�L�n�(�1���:�]��G���_ Q�c��#lݺ�k8�Û4j�G]�߾�wa���[���a�I�������84�lf�;��ІD!��U4�cX�_g���Ep!vn��WAҜ�E�bt���R�W��n/�+p,j��Xh�/���s�����i+��^ ���@Q��+�FjJ_��ia�ʲ�?^�OB�
nǞ"lÊ����ܿ"㲧�& bOG�
�ۑ�����L�[4lXn�)�ߖ��u�	�ժe�.Uxz�]Ã�,�14t��=�����*O@�:Jjue�}�{�QG�s ��X=�]2X�**�Q���_�#`��khf���1qB���9�s��-[[W�X' �:Fy7�ؚ�;*R���0oR�֭�(�u��}\QG�3��Y��]k�e��0r��;�b��/�F�3<rL�T�>~WDYg�/C��I����/r��%�z{*-2i�$#Ѯ�l9I0`��&��E�k���@T�(��۶n�t�BL��j�G5�;6�-,��r��4l���Zp��) ��.ʍ��=�tٲefǗU3�*J����OҚa%5m��<�}�F�C@AS����{L����Pc�Iy�3�<�<��,]�t���@T�(��ٛ�M��-8+#�޸zM��ۓS����7/{�e>�\V�V��d��:�d1��7������0f�8-h�K2W��jU-��5mT�McBbXc�Uq��>�f��' R���$�Y3f��TN���8��a��'�HTRW��}{�۰nL��:#Miд���fox8��]���&j�U�{g�nx#� ��J�rGBYy��f
��`�$��fQq4��Z��)����뜱=�t� ﹊(R��o%=����ZS\LV�ڵ���4��ŋ���QLx�1ʻ9���k��$����oӴi<H��d��ƇNa����*$�'[7m�G�E-��Z}
� �n{&��/��&i�MU]σ!,gHT�(��!��:~b��� ����}(_|��Tc:5=
��᭷�j:���)��?���!���5p9^�a%�M��Z�ȋ5�e�r���hR�q����6N�gG~Aѳ���BwJ���ɒ[��?W�ű|_frjR8��,�t�H�_�@7��˽b�����$��l�ߌs*ګJl$e���5Ä/�6|Q��:�A�h���s�[MzU�ׅ}���>�^''�`��^3���/�l89'��ؔ����
5�F�1>	�(c�G<����_y'�0�C���)QA~y��J|�%	7�i󦛜1wd��Ս���~�8�4k�js�M�&I$=*ry�����k�_�vmR���C�5��1�<��"߯�Q�)�x0�86zP�%	��x���G��H� �Ǝ� �)�Y㋘��%�3���P0�G��Xhu9=��.��wt�������s�v�LQq�(W��nT����KVZڢ�_uNu<��u�� �.�ƗSC3�*�f���|q����������q���{���i�i�R�5,�9f1u�`)zku�y�g�/�c����3ٻ� QƸ�������}e^��E�����P�������0�Q�p��@֬^+�`1֋H�s#nXX�6�JcG��;�p7Ɏ�\t�K�` _\Ѡ���<���or��w��懕�t�.�%���I���P,��>	ȸ��M1;�Q���_`]��x�� � (�Wx���R��6?�{a�-Ikg,*Q\Ć����d�&@�{�I�ʜN��G�����t������cW;�* �L,Rb�3����Q�;�_;G qV�=��B+���?�fA԰b}���>��xV�k�<����t~GO��}�e�/e��ȗ�v�ܛs��~�� A2����E��lU���8"AӰ��+�Y����vʎ�|S�d5i%����ͧ�J�z������ ��9����B�y���y��ҤECI�\�� �b]�h ��/�yłjjIJN3ng�z�Tž��D`н�����qd�[�H^؁��k��Iv���4V���Q#�sG#�b�\Go� ؑ���/��[u<��u���@R+�A�K�B9�H��u����ZUu�5&�����5)�I�6�b�2%F���:�}��&#�v��r�����!&��J Ğ߇*_s�����쫯~��8=�VCu�y\���~�&F��r�!�IjJ=)�G���#X�u��F��Ï<F���I��]h�m��^�W~�	��EoȢ�d��q(I�ǆ��M��J���3Ym�4���" Gr�O>x�=������#:D�  Ve�ߢ���ұ�UVy>g�Ih6�u����'ߋ;%x !7x4\N�3n�^ DO����ƜR�7�P@��&@4�x�Z�TVD��բC���N�~�np!0�Ŀ322H�{`Q$S^ٟ�i�����lx����D���ܷ�����a̟"0�Q!o�'a����2�8i�2$-5S~��0RR��uۖ��g�Krz��
��?�H�&>���[��_��z��$�|�����~4�W��^�8��|���x L~�.ȗǆ="5��$�Ǎ�UhB�ɕ���/�/����{�r������&<F�����x����@4�F����1uJf�,�PR>*��Y!k�M��R#�)�M��#�8F�@�	߳C9�-*��l�_�Հe��L�K\��U��a�bJ D�޲?���s�:kԴ��D�-a6xHV7m�PZ�la�+S�ܘ�s柗[$(^

�H�Y?]���;	#v�+Αe/M��\���"p�_�Ow&O� ^�7x�06n��!\���ط�I8
�r"tW��r`��dGA�t>���Qp�'��Wr~�&>��u���{�����ő�ao��Y���@����r����������b�K���wޑ�~���V��N�W�P��<qvU5� �C4��@�)�T�eh��T��-5��E�3�b�v��F������'�;f�;g<6�?K�� �"c�})Be�7�2��\	bi=n�7��JFl�-��P`�!?���@m�Ĥ^�X�>���o�*���7�lIIK6�#���'M���������1��H�b��h�jMy��J�ƍ���	�*�O?A���^�P��޶ă�S��~#����|!�N�,�~LX��1��9���~w�ܱ���C[�W/ x�o>����bR�z|��P������Z}�+������z�HD���?��ˊ+���Uf��';�q�zJp�~��~��f-����o,%�@��ۿ��o�܄�
0X�v��k�V�a�W���J�L2�uڶ���a+�_�A��yw�HiW�/���o����o�w  ��'N�"^���Q�Mb��3�iIR��$�f9��g� ۩I�Fx�
e�����4�@���F8�=�= s���ѷ1%��`!\f�{�A��D�Y>ot�jTT@x/8f*��'������y*�fOiT�Hd3��{�/o��>'l�Dω�J�7k��  ���mm��(3�>�h�Jx��P�(<�j�P233e�O�a�cr�����w��G#!�����g�R�E�w@���Acmp��%-V(�M%�g����/�M�S�/0n<BL0���`�l���L(p��\�	����?�����KV�L�D�N/�|��i��I߁��1'/��<.�~�����Lh>Å3�(��� ��#o5̿j�-���( T�U�� 4.|�UW	��ҫfN"�T)�b�ى��Y���y`��)�\�zZ'����Y���\�� Q�����{cIvAD:��ϸ���� �[����4��.7F8%5]Z#Wy3��-�w��|�@�� �7^G�+,o=5L��疛�� ��TTj7Z-:}�d�"<�@�lް[b{sD�n�Ԑr�e:,f%�~@�6n n�r<5u�� B��`N���p�~���1t�,��')�Y�2Y��$�����{��[_�}F-�u:��BLj�?��C�0�a%f�0�g ��X��p2�͡�u/�d�aW��~>��ʙ?��g�~6�!#��y�m�V5#�Ǵ��)=�8 %� j�i>퍳����"OZ8����MJk`
�6�Y���@�K=�,�x�S�3 �l��A�э��[���̓%O<*����Yo&Hj���B|�s�1 AP������ ��w!S���/�&�B1�?�8C��F@����[Y��7$Q�N��!�a;Zz��  A``����$�>1���:Od��ƜY�����]@��f�!CM,b����K�4D������kH�rG��ca�i��o����iĵ�+�%>#LY%���^"�G Q0(]\��\�H�)�3�+�{�	���{��{���s�?���lH]d���a�$[�d��M����I;����/>���CDm�>J���?*�h$G���GJ�Fn����L�)�uj���j�8G�>�(�S�8f,у`,���U:�h\|) �	
�\ � �`��'G�t� �� � S X��H Ǥ�4W�<���'�A5���\r�t�֭ �D5��^E"�u�_�Z��v{3	"x�89�g��K���۬�f�um%�w[e�M�f~�ܧn��>̻��IME % �V<"��]y�̷?�� )����6m��o%�%��0�DY#�嘑�w�|F��������  b8Hj�t��VTQ��1�o!T\S��^p��`���� �� .���H��Jl"Ȱ��TnQl�㡻{� 9YL;=�Jwx	*�Ϫ%��RN�,�И0ǞuN�RS;����/�b*��D�H��Uʭ���X��V�(�N0���o��i��9�IU�e�
�i�%�>3��q��:Z܆ ��������'j��!5����c�s������F��Mme����kaj֭[g�j_��qC����{�g��.�O�1��h��믽�
;`�Qt���a���f��{<>H��ɇ1Ǆ��!sa��1��4�{xPQ�i� �yL�<��0D����D����*�1����V�ϟLse�[_b7��AT��\-y%�ҧ�:J|�Ьǌmm CH�i���i�&9�l�@2��r|'���|�*kOq�KU�	&���ĳ(Gq��o���e���W�w�s��Fj����_"��d a��E��MM6��y/y�A�8Lq;�A���0)��p�|<k���pWAoi;j'<�spcc�@ �c %���xP.�AC��
]ڌzif�*\� u���N�I��|ɐG��1���,����UR ا� ��3Ĵ7$uod��c,��:��*�ė�u��a#�b���ӗY�$�Q�����*�ܸqc#������LU�AG����衇��,z�h���:�~҈��|��|����Np����������Vo��T�H�ԗ�w O�C탕�����Ɨ���I �A�2$uR(W>�>VZ�8 �����u�!�0�۶���m�B.�P�Ri����%F]%����h^_\Th5�����8�[�p�!�)9��	{Ճ�ǥW�[<�P���d1������<˽*��k �Jm�@|��&�I����|-|��T	#�3}N���xS?���xi�ћ� �.����6p��N*�j/�T2�ޝ����Im�bJ��*�fV�.�/�����Y�5?$�2��p�z�[��x�B�3H��Ĩ������ �� '�\E����'���5�w~�8��xd��|�P&�A��-�;����T;i��o��jdO}(���4j(�g�][���-v-w"�i�Uq���Z��L��1�5T[ɩ�SD��<.���6���4�F�QV_LMud��Qȗp�G��Y$���D�ke�~�j?ZE�p@�v}�d���o�،,?���m����	�����M(G�<��[��w۶mK�b� ���A�)������K??|�>�ʑ�%i>�q%7������Ŝ����Q����,C�`7�t�C�    IDAT������Iӌ$k;�u�H�'�go�q�2(�|ہY�1��1�-�d��@�7e���C1�w�j2��hۙrG��NL��B+=�wT�>=]>�r�x��D�"���G��f�.���w����-�`��	�`�.�~�Ñŏ�i�-�j�غ�0�8��vB�+?{�����f�$��j�-���	j��>A{8hr��@@ Hp��Ҭ�_�v�QC(��P��83�� D��j�[��&�q�e%�q[��r�����<���3_���hR�쀦Q��!6�/@� �Z��k�5b���� �μ-��F�n����bb��sb�n��&�tW��Rd����;�$����߅��u0�nl���{��4�Vx
����!�X,ɬ�v����\< @ 6Ead]���x��Dq�BZ�����z�K!����˸:�g��p\vXu�]��A� q�A�*MRk�	�4�C\�;�>����	A�����ݝ�n�݃��K`�o���Ч�����AfkvG�kl5ϿKw>3��\(��Ө$�Q��QF$_6���K����?�61w� ��ӑ���;�K��UL��]Ƞvն��O�l�Y���X�f�;���bZP��G�h�bd���^��kv��'��Z�����	"Q]RaS�W@<i���_���*���8�t=}<�H���\����j��&��j�Hq�p��wx�����ϞZ&*�s"f��@�_��OF��p[F Nv��`6T��k��,H������>v��W!��4��Dcl�J�N��]�*`:�޼�cA��/��^���.	�U�����"�?)����uJ��F��GT#��zMxN�������Ue��(Smz=K1�]6����^x�����˳�\����kqV-|���_����r�0�Io�Oprh؈���N�c���^����qk;�R��G�h$�_�&�яi�S��_�/�N�����P� h��r+� ��6]u"	k�_��0}�pC��rL�6sB�ga��a�  8�_�tW�
�h*n�9��ηB��߄@�`�ӯV{�	���+�n���"T��W�X�r�f����2+����so�����n���!��R������hc&��wãH6f�Tٓ�r��.�TQ�=`�7d:�ש�����/k9���X�b7��;�+�ڈ`	��?c�
3x���ix�u�"*ƊW6������B�Ұ���V�g���N+̵;P��@1*�0F�n�ٯ���8\5c�B�!�v�����!0`�[�x�?�A6~����`�]�j0v+ȉ����u��\���@ ��w��m�A
��涉l��l��R�S)�4�� у�Ϡ�D�9�+�M�����'T�^��{������.:�tHm���k9�8��|��X��2*�ϧ1�M{�T�9�8:]Crj���;�����	��R����#8ǃ�$B�n{9�Ү����5F��`���9<-�|�����7�����_�(A�	|��`] f�o�$Bi O�DW��}�c�X4�:	T��tF:����?����.?q�F&�B���TAs�'	Sp�����W�"����s0zIb�Wcn	�~�v�>�`�\����Q;�M/�K�k�U�����}�;Q��'� #5F/�/�����e��`5�����	��*�K8�c�h��yl49^�g�5E����t8m�`LJ�H��  �b")J�eS���$��U��#��~��J+�	����E�uqߒ>�p@���&��[�uh���X�{T��G��!b|c��&&�Z��	�}9���m_\ƣ��w� ���F蚶�� 
�6���V�������i<_�G��D�	˴�ExZt��/e�)=r."�_�_[���H��Ƈ�G�8&�@�[�5������f��uU��fwwEu�R�8�u+��p��9����MA��#�
�K;g@<Z�Ȝ�@S���ʽ��N�(����;*�^�j2�*��)<�Z�qiF��J7P��7n� �=g��ʿ��ӽ� ��&��O��o��@�LeBަ#r������t�u+#O7� ��!f(���sq�&"�x�'���?a:m��=B!�ƨ(J\T���ꊘ���|�i�亜��c��t�T%�}y��^���(|b��0HN��Z'n������%o{Gq��"�
Ɔ��(���|f,��~�ކ֘�e[�[��vg ��_)`9*KW=K!��(/N��NCd�� �
�f��<=|q�D��r�>e�І�tk�W�}G����f�^7�e�\��� )Q`вI��&��ܬ;��,�Џ��b4���>�	|�+Z\�'������?&u��؀�Z(�^Q����4@/��/6��B���t�~�xmI���O&��W�t#��x��GԮS��xZ:�4(Ǚ�i¼cF�í6�``��8�§�gH������:)����a��'�
g�T�������<BŮ�o���8���1g�⼥����+�ğl�U7�Phʎe5���G̪/L	�*��q�@���/�c*uMw�x?��>ˣ�X�q��R|�<<<$�F!7nq�/��z"s�������1@�,} �}�
�E6�C�$g�#�`�GAR�\�imB����h[F�2���Z���b�@�)�̐��BQ�������.|����{GC��fU��e��&�_�i�����2ҿ�6�{���䶕���n9���?�#���b��|_x�,w�Vo���<^8����9I��Z�[%����'`@`6��[@n����u��<�q2+�'R�Ȓ)#w?ܿs�����Ѧ� �Ҳ�}����\w�5S�J�4�5�$��#�F�;�1����CұB�x�#�sڶƷ�6����:�Q��[��[u_��=(v���w���9ã��˿��<��?��_&8_3(�FJ֩�R�Wp�?�^�S&E�G,mͻ�W�M�� X!�La�FB-E�u��^�P\�N���(����������A��b��-��,�*���>uL�V��,�7j���>L�$V��ӥ{��v�P�=M����xWv啣¾x��/��t��T3�I�R���$@�0R���ˏ�_�@&���X������5�hì��<v��+cɾ�y����$�g&���b�����~ТZ��b�GX	�C"��FR����*�7~U��cP+15��:+$'��(��;<���X��!�=%��f���R���u�}R�Y�I���¾^��Z�cJ�B�B���qF ��>b���d�-��6Xa�O�?E��6��%�P���/a�ı��UL��x.��W���������S�S	���%�_�E�-��H7óa��ǯ����;��"�~�u��k���!r�@S�W�R�Z�=41�W���oz�,Ϳ2WD�π��}�b��b�\��}Gp Í  �&�q\;lJ/?��9����Z�w�Q�)�2�IϾ,����i��<6�c�Q�Vg��)ϞD���-<y���	~���c2������lg�J���Є�Ǥ�~�l��jE*{�~'�c��˒M�i���`�l��y"�~ 8���l'�eow�p��T\2��:s��ֵ�? ��G,ĩyxtj3�K�5e�kq��Ղ�Š��|��i��~>�����^yJ��l )��M��[���3���ދ�_�y"��4�,�����1���GG]��7Z<(�a�)���*�5i㨸ǞZ�$��Men��,��T��!3j	mSݓO?��Jܜ�h�l�)jSH�^oc��;5e|3��R����`b�����_i\-M��
F"���i�9��R-\֏5e����R�v�!�`�ff�B-ƽ��r[��4���¨)b����,VU�#�Yy�htGa���Xf�cO��K�!SZ\�Ym���qN	��  ��}ޱ��������N�KJ�,���[���ͮ�G��%���O�����Q�w��h�[Y ��w	G���[���C���vo�n��$S�w�m��=���Q)��5.�����l���GS⸮2�* w��8�-�������V��H�`6	����b�q];Y.���,w�Kдr��;,2`�C
 P){K�V��&P��"	�X��ز媟%# �0'V<54R��@�o�-�D�7C$�ў�JΉCu�HVv�>�#F��Y�ұ���]�֊e��R�	�
r&i�&��5@wP��u{�E!�i;�d�����oZ�0WVH����;�ڟ3���g<w���(ԫ�*
Sil���4��9�����I#��RpQ�Zs]U�z��x>_��c�1JY3��$�g�E�8���D#=u��L;��a�y�n��53�-�i��K&���ɡx�4y����������hӗ���8�~C�oZ����X��ME��m�I[2bXY5�:�uݸ�d���v�4J�'��5)D��A�Y��o)�
�^2v�Q��SY����c���{���:�&��x
)e���3P2<� ��J�
v>�yGj�EUe����:���V'-���D�g>�px�
��A}����4o��|f$S��""��D�Af��x-������K}�>�k�w����������P���:?��,��} =ehʫ�9; �]S�V�,�_7��l�$���=��.�+��Mu*���{W���G�6$����%t��{�:����3�~�� ��(��"��,�� R�#�6���_/���\%Bc�]��g����^�޸t�����J(�A-[3�&]ʒ��h12��Q�t�M�Y�bq�|'$�d��V'���G�~��5g�/'�F�����J1e���,��Ÿw3
�}���9��ׂ4��������f8��v�Kٝg��,�T/�ԍW
����۳��/�a`�3�b3���٘;��%�	�u���U��0w�6ݽ�6.����o@��=>,\�F���ka�*���Iq�ȶܠ�a�.��z�@�_�[u	�:7�jB��a�/Cܦ�%'�)�t>�������SH ?�T���XS��n���
y/�pl~;�R|�J��O('�|�5�z�S�?��_��(2�0p��p��gA���'R��Y�������m9k�H��b�;}��>4����4y�j��N���K�	�"\��<���D�d��E?�a��cj�b��鶭���n��?V�����\i��"��L������qU6B���%1Z���O�<%�JS!$N!�w5;	.O_��4d�H��A�{tW**���7X�(
��W95�>��=��*u�Y���Srf�o�����R�Ø`@�5��|�}/�(���FWka����_C�0�ى}�D'OA���'����6�E��2 �k�#���1I�k�z����la��M�p��p���,׷y�����$=�&G,�x/�v2ξWͱ7}�2:�H�%�{��B�T�<���7L2Τ6�,{}mp�P�r�]U�d���H�Ȑ-1��4���4Mn8�(/헣�f��*Ҥ4��D|��9dd�	�����O����	�6��?��/��iw���Posj@ai��B�h�ΔSz0��ro����ҿ_a*:+�;�'�e�� *� ���$)HڛTā���x�b"�P��H_�d����I_��G'si ��57a ��ϵ߯YF�G J�RD�zwsx���Z�"��(ὅ�|�}w�g��,��ē��I��srd���Q�V<�x���ة{�E#��K���J�Ճ Q�V	��U%��u Kl����{Th�cL��@�R ����:��K(�A�T�P���-r�U���F��X�֐d�VJV�x\2N(B��s�'�%��k��6��7�&�iK��/~�U��Uj�;
�����&ן��ō�����~I�r�l����v�*T�OG�CGF����&<,�>������%F ��^��,���$�4� �����e�8���ډEXUw45�����8�@�dp��华���TB)�s"� j��BҖ�%2J��$�?��\�a��n�#@��p=�̊~6	�=1g�cI(��@N�P~ 0%"��x��s4 ���.�
�"R�b�Ϸz`D�W��ahK��jڂk �ˉŴӝ� �k?�t?}��Q%F�f���Ӥ�I�������ֈ.�Wd;;�Yj�Tq?˾��(�3�)�hѵ�E�.�L���>�Ǹ�?�iSi���˯oW�lI�����
�s�2�@f�m�'y@��GH�U�$�	YG��A�7�Q���Yo������J��$�I�O}9�3	쩻-��)/� ^EJ�G���l@�H��a������&tP����<TD�����O`�T*!['���m��?S	'�ʑ������Aك#)}�l����E���^��@,'m@`I:� `�����kG ߄q,����i7N��$5Re��y����:�'��[�̜�S��(C���.�ջ�x��Ϸ��`t�W�6�o��I6���'��^���CB��tbw|x{�-u���O;��"8�X�E�

�"�;AU("3cf/B���m;�jqMe���9�k�AU����bo�������fj0��W����Q�t9٤bZh�~1
�T^����. d���o�-r�u�yݟ!cFq��$�" �h+��J5������B�ra�w���N$C�PgKݶj`a��ʥ����oI�[�P(�+�=��?��%����J���n����d�v)	�^Ar����I�`_㮼�nq�O�|��$I� �gER�N8o\.݀O����x�u��\>��
��r��E$��c��V�C�jx9����߉r���r'���_@��pE���oOdO�)�����͝���74��g�!K&��!D�'d+ސ%��@hL�Jգ��t�P�o���
�����dI�·2|��"�oXA']/B���-��Ͼ8 �O|b9��$��S&&����^`����\aX�D�H:~��4J��=��518�e��6e�
��lF�-.#�3������7�d�.;�TaJ-��hT8	x�� ��ៜN>�AC7��>a�ؘȜ�N�K|���חO��MٴBҟ��g,%�:"*?���w,��f�,.&�����;�&UP��D'԰g�)��n���eݿ�^&�{�]Š�����|�R�3Yv���6@�X$,�R��Ϋ�ị�n7pB8���� zq^��?�#�oHO���P"�~6��>O���&J��M��G]�6�	������ㆹ������
{mX���/��	|�vB(�8�e�S�EH���=-W��r݃�wR[���9��b@��bH�>��YE_mL��.���V�3ޥ%�E�V�Yb�u��oj1v����1�%��?cg��?eZJ^|�*Qf��(,��S��j{;���-�����jt���륽�I����B� PS����/�ªWS���.�nRughr��o`d��֮���Rȴ9��xy�TS#
Ψ_R�k?n9�X�ݗ�}�iST
Q����/i�S��ߘ�R��)\6&��?��ىc�|_�O����%�z��ZJ(ۺBu#�_"����}ظ�)��5��Ց�q�ΐ��c��v�Ks�e>���Zi�zzś-�~WI���+�4��I�ٰ7@�i��w	Ns)i#�2߅���6��,�]��D���햙�ѽ�s���HܕDe���Қ��T��bɷ�i7~��W�&�_���	Ŵ��:�;�,����M5ds)S*���rE^{�_S$Y.�p���/��b4���:�ʫ|���'M���rl#�f��Kp��=��>D�)�]/������ʈ�&SNN��V���֥"�L`���%��)R�A� ���z�<��9���Ͷ��&i�U�Sjk_"M�t�a�p�@=F)�z:�R	i.5�S�=����>Np��$��U�J*Xqq
w�����e���n*[
�/jjx����)sMd�!�n��!֖yw�Wƞ&�_�?n���4á?������^�@pn��A��=�u%&�Ve���#����Pz��ِ�T×���֡�ɸ�r�(�s�Ϥ�ί��,�>��Uk���0ܔ3W�f�,ڼ,[�3%�^�[細"<��J�f(�#՚��$����uʱI�Xb�X���\[[ʴͣ�>��s޲�����am���S���^��T!}d�K�upxQ���L4PKT���$�i��<���"! n��N]&		��w�+�;��۝�J�<��W�|#!G��A�4Z��֍�����5%��'l/���oI[�KzZ��5�Ĥ1�I;y�]��|�����>ʪm���@�h�}G�)[�!G}0�� r������K�2 [������q��5�����%3'LvR3s"�Ϛ��38�WD@��#�˘Y��7�i�X2ISÜ="���Ӎ��$Ot���������o����0QŤ����&�7Y�@`p��̏Geo�d2�������q~/��I�@�ii������Sv+m��@���@T-�c���rX�I"�~1� 	�΃����AiK��"3���b�,-�&�����T6������^	��ǂ�u�K��{R�	���a�,���J���Lۋ5S��A\��s8M~6C�N�'�g�<q>*;w����7���p�&2�G�9���?�����z�;�ʣ�����.��f�����h���sM��m�_� 
P��`=q���k���e�����'n�e\��8�;0!!�@`�����e�y������ګj�c4j�w�JK��m`�����b*�y0�ܰ�5�L4y6%��-��Hj�g�e9�/������m� X�����=`�酩hKZ���/�O�����?pZm@7<ny\"%������4K(���l��5d�w���U���!����!�_~��kg.N�/f�����lA�,y����"NŬ�/{tU��©�q����`������t�kxެ�����W���9= ��仗ٟ��ף�% i����\��_�L�������!
�5d�>r~g��z�Č��
�,�I0�Ww�)��T-�բp`X �m �DD�#���W�9P�#��ǽ�ÃH�Eg.�D�2��I�����9;ޑ��w
gxawZ �5�zx�`~�aӵ+�pM6�^Q��4�����{��q��FA<,D��"�&P�J_(j'�6w|wk����Ի��*��ʇd��W�i�?���l�b,���Q$8p�v����°.m4���UF"$D����T�
����";5Tp �@z��3���φ�"\����E�L�j7s{c,z��
(�!�K�����T��,�b��&d Y�ӢM�rz,+�#V+���:��2@��������g5���v(�`���Oe砙$ oAh�[��Lv���(���(dR+�ſ/]��k�N8�'�rm�� �a�8�<�Z��hT+�x��5':E�mQ��=,��B�4��:0�a}��J I�MEA(���I���B\.Z/�5�tp`IE��6��G����4[�^�6u���T��;72�:n^�`9�ͪ��`���b��Pq/�w��i<�n��^�iHc+h��OZ���5a�z&��͎
L`<�a�ai���")�hBY�sl>��ús��8���0	?�.�X̕*o����gEY�?7f+�ۢ�6�BJ��-�,�M�}�I�K�"��R$�a���=�z{�5O���u�R>��$3Y�-[��	�,�� �}n-���~�wI@\<��������fcM�lpP6��p��̉Γׄ+�	�|G\18��	B�7�e",���'�r�4������5j�.��K���Pg`S�b��h|pW�����d�a]�JGC[A�yCQ5�0˸��]	<\��s F��P}g|�e9�1J$����#��\�A
������<���>�u��dt���.�\�@l g�縢�;��;�a���8����l���q�pŁ��@��9��F�#fi3�)koG�<�-���b��j�~�
?h�IB�A��i �����\sHzy���H�y�lI�z��ǌ�7�9�Y=lm�篫� 2ؘ2�>�|}^�0 �f�衉��*xD��� a���1V#�{��������L���@�ڬ�c.�:�ͧH��&
�52O��B �ҝ�
��s s �ױw�~��� -�뎑��^,�����SS
Y`r�}
r-�p�E&E�{G��Ѹz
�_����(>0��U�~���er��z������T�ň3�����]�^b����o8��0Z��R�G'$q�C���K�[�y�b�t�6%I%7V��Te�d��P����Ȝ�>��0��3u����l�Q���e�B�;7~3� q�'ԉx0+�vK�+0t����a~�(���Bʻ�g�������(%L{a0y˻ Z7)d8��}�W�/}��:y�_c]���7^��(pKt<�RXYR���\�gk���`zwq��$K)"Y����8���_�*����/)�l)�d*=F����;a�����hTl�B��M����qML`2y�����.SK�hO����|��/�~��),o����R_�{+!���KU:�p�e����u)��;�~k8dV�,L�("�+��?q.,^�Չ:�?��V���E�z��W}������^q���Qê�]�ƨ{�'���t��Ҙ�Q�
��,pZH�a�Ft����RY�������	��vTl@i͍=)WVEր+��z�"1�Jᐔi�=m��L$����)_�_煁~0��\Du�5�A@a{���������茌���`�3KƓ6�av�KOx<v���[c�����t�鞰�.Y��m�
����3���B�CC������
^�"����-(�$�80��*��晏�(`k�8Ջ̭��N�G�(��#���B28���u(� G��K����p�P��5�j�P��=��ÕU��)4R��p�8`�L8�S>+��W!�O0Z)uY
���V>0k)+�����/�������a�+�^�}�� �I@T��z��[��g��e����	�딫����~ yCF�c��;�)�r��=�$�%$�q�B���!���IaUi�ql촰�]�a���8�}��.�*؛�8��*��AӍq��#��������TiF�e�Li	�yW���S�w��KPZ_�rM	�b�tW^կY�+Ɖ��X�!����gL��-�#)h���+x�7�W[�yC��1�-3��g=W��f�Q��61�eJ9
�Yj)7��:�$^߁�P���z0����!���;Љ�P�ʏb�,�E�31G
��<�L\�a�6+k�_�+&�έ��5����F��`�Ao,�0��,%�U�v��fv�zk�̇`�>�?$��j9BvѮ�T�r6݁lêϟւ.�Ĩ��Rgn���>P#�?�/>9�htk^Wgv�z����J����hL�*j���6�"t2��x.v�k��o�&Ic_�E$�n�oB�N�l����y��ST;ѝ�	���.���>��|�3�TǓ��Wc�o�w�G�Q����{����C-6:���.����D.�K�U)]���Ovb/V��<v��j,�����#?`�tyG� Ѐ��p
C,������1X� �\P��]����?�C�'�l���6İB�n�6��8&�-(�IX�
�����_5#:��+{�_��!<����1������u��aL�d@�7��ɍ�A�L�	932�ێ�[�T"6��׫���_�vC��K%���6���υߕ����]�EpS@�20��\���D�������V;�M<͔����G$�����Qc�;��ur�j=��׮��՗�W��&�O��#���tYSk�I�1��\Ռ�\�!�5nۮy��	-*��F�M�u#�����m!�-mMOR@p����<F@���E��@2۔~EI�����9�O���2����ܿ[
�X�`�)$���N
��ʳ�럳Ls��^^�^�+Q�8������[d���SK�w:<�Z5�bT��h����$��l**,k�'�P����ބF�Q�H�vc����6%��4�j�W$��][�����X2��^\��� ��u�����x���[��$n�v���M�@?���4�CbpVi$�/��=�X�Hč�O$�Pl,|�XU5�al�r:>"(	�'ʈ�q��ma��*E6�2�V�Oת�cfغ$� �!Ś�f��O���m����@Ll�'���3�^@���J��+��WQ��� 0H[�-�!�ÑV׫~�;�~�����gz����f�6)�	}��gU �%C��p�d�K�k���ӟ�G<>�*�*�L�������%��\���a���1A�^��1Q3�%���c��3����~i����l�H�Z��S�;���\��xI?�R��LT�����7�HH֚�O�!�Ϙdox�����&/\�f���g�Z����(�J���P�rMNS���{�y�B�^�8�2�^t��n��J%kwG8 �oT=��	��A)�]����q��T�lѓ��(BV3��N$-��������'�:���!�n0���.+Å>�_�9)�D,xC�T��\�V�]��#�=G�����c�iM����v�Vt�,,��󉅺��9Ǿ[���H��%���-��M��R��j��B��v칌���.�H�<է�FS�z>�k�F����v�
���F?K��|�]�*	�V��y��Gn�.J^��+s�w�G�]5HCe[����#����XW�e�H.G$�-u@��q����A��y��mL��MdcQ�a3$�,+u��	>A��f��'�;~k:��T��(ݢ��8�99�D��%~&�eJ<��f��>��v��oSEu�z�����L�oJ���<�RSk�p>�u�3��r��/�{
��ӶC~Ɯ� ^v���Ն���uv�:�$�|Q����`��/�b޹��\�������K%��g�"�p|�#��|��j��n���?X-�⿲ߍX]A��S��gW�K0�Y>w5��s���ƚs���8b��6"g�n�(�´U��T��0��q|G7���z�נ�r?"�*��T4�X�"��jF���o�� ����'V�ڏY��É�s?Qg���J��5W$��Y�	:*�(,�6����:�x�4eO��U����	���}�K�<�l���n��ih2��Ў��ps<Cs�Z��馛��*�"��E������ޗ��'r}�$��j�p�ɭ��;�}����;�UM��9E�-{�F0M���2�=��! ]�yI������5�8\p���s��X)��Ml#��a�B��:҇�I�W��*�W�AFA�� �p��U���A�_�(R"�<��S�T�� ��Rm�3��� ���dT�G��Eep�eTD�ApC�4\8�����x����zO�v���3��+ȃ��O���M���PL�0M|��-u?i2&$��~a�~����C�{���	0�z��;RW���7��o!��z���e�󿏑��'�.K#�U�Ŗ������ �"�pG	�K����ſ�)`�4^'�ÌA����O!���+_�jQ	N��������i܄$��(�@	f�ݶ�,�f���"
���R�!p\,R�澯��V޷�|����L�4�/�^kPI��ǭ���aU.�6M�2,��.Ug��)�uKB�])�ً�c�j3
�)��OѤ�.Gʔ\&l�� ɔ�0����M.����r��!�u�Ѵs�ь�_i��Mi$OՏ��&µ�e&��ᰙ��ޖ��|�M�RЏ��kdSe��m�m����]{����dX)G����u'0�f6�4�P^A��K@}We߸�8jyVk+,�+��ʑ�tʉ�#y}yK����`+,�_ŗ��C<�K������;��e�f]��Y<-|�6�m�8Ñ�lޞ{�����<c0� `���J�7�
�	n&�M���x�||�~ÀW���(O��1Ͽ���S�,���d����E\y<��s�>8�6=����Ӄ|йA_ft���H.AH��)��ê3��Gg�4o1ڢ���2a�gߋy����{> �@G�/���`;� C*[h�A�f7�2�D��B*����L8ֽԢ#��?���>� 3�S���Э��ɼ�#.��$����XY���}Gq�wf��p�����r��&sw� (d�W+�f2��)���'36u�zꫧ�Q6*�I���\V�1W��ɕ�6��4�J���މ��u�]L8d� %�x���o�M_�<������ÿ�Dca�|xƢ ��b?�yl�:�j�䒊�\i�<�ơ П�N�xk��X)D%4u'8`��JG��"[�ru��~*M�{�P�,g� y���N�s1���6�\� ����.���cΓ�}�rE����1;G�=�z!��a'ӡn��֕V���f|��@��\f�%�aՓ�a.���D�Jpk�ǔp��V�{��[���ږ�(���ʋ���P���-��(���`��:6�X+��ך�I Ly���7{{�al��V���#�Gf����V�K+��Jb�B҄  ���n+@aU�[�X)	Z��m���*�O
@�%s<6��A�^�* l�_I�\�@���Dx�@R"$X�X]���i_v:x�.�!�Y����S����^lT\Zr�����	O��}��Zyw����!��#�ڥ���u���&p����8[�F�n��WH��I�ZַK&�1���><��4�_�S�cl5��Ϻ��A�5T��a�m���nǳ������)��lW:��Y8��3�T��1Ϙ/�Y�msBK��x܄>����U����cp9|Z�`�.6�1��p�cڤ�c����a 0���u>>�!���2l�k�?���[�֬8�,�
���*2�����XtK&���~���W�T��;�l�MG$���!������EP 7�T�t�m(��t�cqH�q��i�n�/`�I}�)f.^­Dq��y����hu����'���������u7�i&��*���<{�Bw�`ʷ�����'��^����ʬdC�2��J�;k�X�0�O9���
�	�`BD�
�P���Z��� m��}��-O��Y�&���9<�����ѱ�	b����_�-y�3�Zѕ'ʕ�>����G\�r�V㽯�Y�V��d�)f��xNxzzm7~���G�%ѡV�0�����%V�#�D��%�:��7�Z��������Jv�S����� ���l�X	0����͖��a���I�2�8�Ue.X���	�αuM�%����L�΅�I�7�ԇb��2�f��~���κ�����AF�"<:���_zӳ}M��fّ bA�;�ۖ?l�Z�Z�B�!��=������X#�ÿ���8<
�^ei ��*w˴��?	�a "/[,.�cIUah
�E�����ߏ���3��=C�|<��<��غ�� �d��#K���mn�H� m�=r��7g��9&ߓ�2����J���ۤ�]����[V�,C���~�z���2t8�Z�����{7��{+,����a1o�':m �q9���@Ƞ{�H���5A�~QXox�r��������e"*��̵�LJ���U���*����Ј��Ԩ.��d��FjʪĴN!��S��vNf�I%�R����Z~�:�fiq4�W=8�f���ƴ<D<(=�"�i+CA���:���n���y�f�b���b��9�S�'�	}	I��Q$幭���)�F�3A��YĢ���z����_|BE�8���Ҡ0!�0�R��0pck�֠5�R&�}�Tn�wҊ֬�|z�{UN��!�e��)�`܍�-�x_܀�Q��w������܎�cF�����G�(�����y'��Mwj������y������[����S���gK�j�~�]>��&9+���O�T�C��mx¿#�V��(���{7��������N�/y0M*G^����1�6@�%2�&*��T+n�b��6�������*�s�a��V�ܤ�� �F�U��$�w��5@�QfQ��q�(8�𽦭�`i�ޘVM��y�#���w����BT���&{���b��~��@���fKtCC���ÁR� �BX8w�NT�|uӕ�s��1�!h���({�޹��bA����F�44j�)�@^D�P)�O�o�}޴IeL�:��Ry6H4�Ny*���D2~83����8�!���'$ǝ�.(�U�>v������M�,wŸ��$}N�8~�����Ig�w����䜤�����Z�Γ�T�*j��|7�F����d�򧋫�
`څ�o��)�і�D-ä��Hp���8�-��xI�Bz�3�n���~~��W����^;n^���l�z�y1�2���;��笽��%� �/)ll�g��-���&��/A\Z<6�肀)��]��TFt��x@���ʶ���A$*�k���x��#�m��A� H���å��0���)Y�5^���ׇ�	Ap�`��I(��:�nT���H@�~Ȓ��]*��4p*�� ���� 6�ų��u�9rx�yj�u���"`1��1��6o�]֬[,�H��ͤ�~��mX ���l���M�VG�]�3@\�6mX��6�[�o�)9�o��_.�Hs��̔bp����������<@(MYx
�yw���swח��b#���܋>WJmP�I�Oh1Ul�+uk ^@�M��Ou�P.���qB�C�!
���󠢹��5=��b��d�D(l�27�n��Ҿ}Vx�3rU�K��.�bO��b��b�d�pz���� ,I/HiW�fz�r�A�$J�>�S��-�~���H���+
q�v�l��_z#TW�  �P��^篫7�Y���#�����[���c� +�_!7�5u!���29$��_�BC 
Jm4�ąU�_5�4��]��R�����h� m�}�Y�S j��>sI�Q3��JjJtC�XV��:&�y"��׻0��@����Jd4
"���^����&?��p8 �g'5��'��B9�
фmF��T/�	 5��\,Q=��XxG�x�� *#�"�i��ET��Cw�U��:�Q:|��BG��/�>ΖQS�KS��XI�q�vi֢���5k� @�u5����m��~x���_�jބ:�QN� >��S��J�jv=;ꨣ��/6�V�.D����G<qJ�d�Yr�2Mo��㡈��L���QKnO� 1� a�bJ�\��%/c��>'�^�0�H���9X�ج���F�����f<6a��F\�����hFKiy�������ٳ �IN����qj#Bio3o��E`F�f�Sr�����`����U*���� [�sp�h_��.MZ�'��Y��'<�Rɨ� �lb�~l�z��� 3�&�dȄ#��5�����B��gHZ$�-G9��8F1 ��v�i�7��)�� ��w��E�v�Tj��R�o����`�� j���0�4�!& �a�P^��8B� �`��$�ʫ�eUW�d�_�E�*L�ƅ0VP�s������D�$���;�,��3��Y�  \>�����`�h|�<&܎�`���όW�&"\�����_'�?Nl��ϛ��x�qV�d�h�W��ր|��-���Q��d�vm${{�lX�W���Î<R���F�;�TY���{�U�}�g&�R�л��=۳����T��ҤX�bWZBBS��A��� �*zW��Cz2���:3'��x0�q���K&3��=��u�^{���у�kq74�Ry)))�N�0�S��+CK�,ჺn�:����:t�6mڔ��(�P��%�Ň�������PYg%�+� � �3p� �� �=��pH�ޭҵ���;�#������A��{�����xp�ԥ��2jq�9��K}atݲt�R�0e2D�@�{Dn��&����S��0��M%�"�Y�`E�[\�p?Jm�x?$1(w�W��Eo�I�����x4h��EҸQ�ԫYzJA9~� @'��"�"g�1�H�y�V�S��ԨQOy.��ueێ���� �[I} XHǎtvqJsqb}� "ۊ�B��ڵk'=�P��Ft�ށ?yt�͉j���$u�,�?y�O�n���bI���q�J��w���}v�2`�pY���[�F?��\M\=���cY�y�?�"R>Y��W2�Ù �y��C���Kapc��Y��8�� .F�0������ 	p%��`Q�� J<:0(�q@>���U�1Vx=�"|�!f�Ӷ��\�zg��KG���j�K��֟�!�����j��l+��P֛t���'zR�B ��ۯ�29���U.�4��>�ө����߫�A� &�آE5碩���������C����\���7�C�Q�M���@�����`���0�C�N����[o���/�*���F��ou�5����v]^�<4����2��#�@�2�˯e����6��cm�m������i�v�1v��fMRZ���	���ju`�C��l9
`0�����>R�6�X�$�K^N��a��lrc�k�Yc�^��ʻ�D������R2A<^E�z[�z>�wV���F��א�F>��J ��
�[�C�i��4-r^�F��_
� F�aP���n*Ow�YL,�K G���S����-H#I�(���⟲�N�`X���ړ`��A���Q��@3"T(�p�I;V�V�6���}�� HX��.[!��C��}�IӺ5Ќ��<֣�� u�s�ʰnm�q�쯾�13>AJi��x���*�#s���uLeB��D"%�H=&�Q���>��+�B�JR��&��dW�1����܄�b;rJf9rD�����4W���:*Ǐ��|�<�se��tW�~���U!-��Y�(�)B/dn��������ì�P��J��\�����+��7�T+���__���[�uu�!�J29������S\9��9�C5j������1�E���2}q��)�e �����`er���w�-�].�/��I�u�rU���W;J��U%�a�����\����&�ޣ�Бm��ʤ�?TT���i-�\w�m�<?l���3zU3ԃ��*�އR�D���V �|RL��5�X�\5)��" $4 �W�VMx���ʕ�C�e���R�^=5��jAF�Z�e�ϻ$7ω�>dJ�  � ~��>������AD����_7+���n}��+�	P�@3��{\����]��?�C-%%%����U����}�0�45W|��M���͋2l���0@�ȫ�#�a��6������֛�R]�^�"[ve��%��SrF��R�IǞ/K!�yg5�!�C��[>Y�J&�Y�x�<zߝr�5g+��~�f˚����jX�� �6(�a��"A��� 9�*lz!�ڧx�jժA�5ރ[b�F\יg6�?o�Ć�3j,PE�c�/�����S� �!Y��$�ע�G�_��)��8GvYo�Ps^d2��A���usR��<[i������[�A�|�	��\���<�,�	����R��o6���N��1E�,G�T��LyE��2	,*~�8|�{n�{�N��-�- �c����Ҭa])B,��g� �U���T���/V�3���ڥ�����_��~@z��/[�W�R#C<���7 ��nd1!ܤj%~�\_	@�2f/����9&{v��u� �������*'��F�VP�C�3� C��u�;�p��{�HӅS�Cokr�eb�,y7d6B �4Wx/�FV�w����k�]�cv:N��M������+����ن�D�8�`�t\_�����N���ϹF����:K}aݨ*b� �1ma��Se!������	����/:WZ�DFV�/�CG�$q��wݨ~��&y�,	��F����MW�^�-k��,߯ߪ�T/���\z�G��f.�Z�:B:,LaP0��!�.�]昽�!WͰ��jV��+ŐϨ�0SA^6@��ԯ_W�n�&9y!�ƾI���f�:���?*�"HuXz4n{�lE�l~��DT�m��G�	�Abj �����U�vj��~hYI�ꫯ�1Ф��<�(@T����_��{�χ:�a�ȑҴiӓ5�r�9�
 �.�,Bes ���vҋ�"�cE�� 2}� ��Q_`�2��dԻ��
�� h�c�����	��3��	Cm ٭�?V�F�o�D����3�9��BL�	��I0`��x\Q셍�&�A�_�cQ�� LYr��kժٌ���k��%�A9o7���t��*���1)*	Ī��G�,'#
��8~ ބ�(?~ �'f�{���J�Q�4��Z9z`��Ő _kO�<�j���;��DAA�lٲ�$Օ�&R����Ϗf1U����qe�G�){%P�H�W`�ﱏ9
+�bP3A%W#
����� �ԂБ֗:K1�Ȋp��9q3��a�����$/�L�;�$5 ��B(��K�&�
����>�i3�V��lڴAU<_x�Ūo����6B� a�CF5��1�i�E�ʏ\k����M1Ԗp��P����(� � @� Y��5�� ��g;�[�,40hrZ�$�P G���3'��o������^(Y|�?^6l� ���3�? ԪF� #��3�|�� /��	]wq�6�a#R/�V�2'�RE�kP@�rK<?V�l�S�L$�*��g�'XQj��oHw���c��Ǉ�W�^Tk�x�jy�8�����= 
��8�9���q�F�����B9��֬�|�/������6�=	������ۨ2� � D��p�b���K����h�$�A�\}ε�FR���l'� ��U�:�Ti�|��P\!�/�-[��;�լY���H��.����O|"@PrɌl"s,b�T9e�������8 �*�aǶ B?�3 �� ��AW�l�4��W�� �=Nt���!q��s4������ �9�{���G��ٵ�g�(�$�5i����~�f7V\n2��s�0#�72G?�&D�X(��Rz��A��fa}<�p�T�9 BN6��hd�8�����$��8-y���ZTMsB��D�F���PH���%����ÕZ0�?����#Hs�S�Ms-�.gN��Ǡɟe����~�Q�a�o%�Čp������tK��X	+xZ�1� c�P�/���EʉX>� ��50�3p�,&(����A'���0�(xVa�����Z�F��ܽK
�U�~c��|�c��~(�Z�)\ �=Jj�� ��lZ�� L�`JTGL~z" �b
�BR�X����N=A<���T}���a��hX������+R?�,��\��a�����=�8���E~���ɓ'#٤��¥ �Q D�Q�(�.� t�+CEV���0� o���A\����u�\��!?�z��H���x8alUfb���!"?���!|`1���KV�{� N9o�je��� ���9�զ-�NJ�"�K�K�q�����0/@x�+1����Lsu�"���!�~�	91�Hse�T#�t��کr���J�!����hho��_����q2��4h�޽�~�zu_�`GEY]c�<���o����H���ߨ�>�aÆZeq'� Q�]:R3Su��1`)M��P(� ������^y
%�ԥ�G,I3�^�8��0�^p
8P��Za�X-6"�=4s��. ��$�.��|�$X�`�� ba�2�Z�v=�u@�Z��`��_�zN�>(qpY��n+�Մ��C��?`�� �鱘��Y�F�	���O�Ȕ9�!��@ )ί�J�? b�? t��ʕ+�w�Q! D��(U���EyEn��8����{��'u �fYܙ(@��AL[�+u��tSO�0���b@辛��ٱUVoZ����$�t�j	I
��� ��Vd2!<T���1X�[Qa�٥ 1l-����.8�n�>&Ͼ�&��ݏp��&��a�9q�+TK�"��r��!��֑fg�	��}r``�p�ŭ�מ��� Jv�1),��� fGẸ1lE�c��& pp���*�� x=F3+�Q7qf���k�'���F�8L��0��7�ʨ� �A�� +�{����^��c*�5z��yTb=}���^�رc�4�I侣 Q��!m� �O v��x�@���!�q��Qi2g��l�B���+��ՈJj���nB30���C���yHo3�oA-5X�0.��
��W
^���2��we��]{دP�V���,����P�B�X�U�;*�6oQ+�3�<G<�Bx*��P5A:<��0X�9���"Fe�={w�2p!b�W H��N8 fK�ԭ��SK,� �oؤ�ys����,R[Q�&��9�DHld1 �Vz���|���(�.r:�u��s�F����Z�j��OZ^�u����R*�� Q�Þ6��^C ���0�E1��E�ܸ�2w�dY��J�L$5@�:���.R@���1c
�fS,�C�M/�PfΙ�cZeǮ��f�(I�L��@�_�Q�����LW=��O۷�O(P�]�ԗ�;w!u�oIR�J��� 	P���^�W^~CZ��X��+4�|�Hzw�
�T�-,򧮑���!ҫ�+�����Їs>��_�<��5i�p	� ��Ȱ�R#���ADJvS�/55U�;|p���At�ށ?{�=جK��8��A��ZϿ侣ğ��c� D���Ő�檛��q��|9�5�b�<�b��A��E�x��>G��TR�tt��l4Yaf� (��<�����}Gd��I�>n��|�z��:�JL��s�I~v�lް$3�U����4�
? �Rܐ�  �Οݴ���"�^O��ր�|�1	��]�L�u��%����ە\Ai�}���� �%NF�?Q���Iϗ_��<'.�ґ����i��΢���&���]Q�QIMן���͎r�b�Н�N���w�,���}W�ѭ�ס�i�qZ҅^�#�H^�j�$����qx۶mQ5��R�I͇�_�{\`�'�,3>'?~�JF����`�l���K@>�U�Elܼ\sظ��vN��`�ep��䏖H��zJ��	���}���,���Ңy3ٴqV�>�-B�:Z�l���lD�4BE,ʻ���{�.��&g�N�������bY��3�ҥ�:o����F1���+�P���8��1��K^V�<�by�gx(�f+9p^�\X� �+������b���DI��	V��kG�[�� �L|�cM��1c�H�ƍC�8�O��-W]u��E��:�z�P�_�EI�Rn0���`WDM��x����d���2e���n�I��4�f��U� ���(������&`��IC�(�*�����En���4C�����2BD�zg�U~�1ivF#��vY� A�U�$8�
�rPY�|G3�0x��ty�Iiլ��}���@Bcѧ�����D|�Pk��X��G%8sn_������xj�����}�Wޔ{:=p���Aԏqn�;4�/��ez��<��2�O�>�)�G}T�����R�=ڟ�Lǫ2��ࠋ�tM���ի+��:�g�馛nR��+��!(���(@�r�~���a�>�9�A�ж��j&�"�Ν%K�,�Qi�lC��K/��x!�a���bb}A���!<�e���i֬Yj%�YI��/��Ͽ,}�I�� �9�b��}r���Y���٬	�=bd���;	�uM���p<+~@�otf?i{�c� ΐ�w��X�,�\�N!�AY16��f���g��_�>�&j�}    IDAT���r���R�[ ]�{I�v$u d; �� �]����� �	i>�$�b�C��ۏ��H�Vb���_o���g���.:���CJ999%��8�~���[�ׅ7����w�D)w9 �6�S {$��?+T����̛1U(�ܰQ}ID���>s�g+�#0{�ЬǊAg(��w�bb�C$�C��)*ȕ��Ce��ʡ�"d2Pu	,��(8�]v��� �W�$t3�D42 ��~�d��_���A�q=M���<^KVVK�� ��;�B(͕���d�!zS��ՄJ�}���uy��s�0�k��,k@��I�t$�h1��?~4<�,&iY�Z8�P�څ$	�ѣG�����\�|��� ��t�{�D���+�Ѫ�ы�>��;ռ�R7���x��dϞ=����oݺu���D�$ 1t�'C�A�b�O��IV�ՍLyK���J���Ge���qM&3��ۨ�Q����$42����ߌŨЕ�I6��MU2�,���_+9�8����P�A�m9z$�}�8�Z*�U��.��N��j�z�dȠ>�2x�:��L��B�	CdP��l]��!0��a4��R�6$<��a��X�6�H�_� "�-��5sFW)�IZV�( �VǏuC)P����W�^��J��ᦲ���y
���=�!&����W��X�1c���*kI*Q�<�=mƲ��'�Ks���BZ)��7��n��R����PW-Q��TE(I��K��C�P%.a��F8�~�?af�h���g��_dޢe�{��. H4A�Pj���u�d�d��@&��1���aB!��rq6�.��O�UI�DB���c3$N�[��!�Y��#�B)Q�%�� �pl�	F��
Ry��	3�(���gO
�=D�/o���)�<[i ���0Zf1�!�CK�	 ���� Qy�@��%�/q°3���J��o��n�0(lwKY�����|�A㲸بQ�]N�� 1?�i�\���9����V�yaR���AʩRh�F�犜�)��)	�؇�M!�fg4QqF���H~�� M��.�̓����V=Y�h���*�	�?����΃.�<�b�ŭ�+�yi�M*}.�-��q!<�����_J����aCx���8(�l��$�]�ꉍ:��N�Փ�~��je1I����Vm�o�rT�c%��S���!����q|j��N��[Cvօr�?�ǰ���i;�͞=;b*�)@�H@0�DpPM|��dFv��V'B=6�$�PC�~�jH�f&�:K.��`�Y�� ��͛7b� &��Ȭ��R,�3�i��?[��T���RlB�$��à�8ۇ*m%�6C�d:����Ŀ�a����d
��3P�	"PH[e��:h^D'H0)��8JI�Uj ��@���ΓPkQ3Ɲ�nְ����⼨^9a���{ ��_-o���:u������1��A��^hԮ][���=�s���\���<�:�zeq��D)wy�EϧNY�Z-&�o{�Ί�0�.TT����/�h�i��]K��0N��G8�k��IҤq#���N���k}6:v�"�/��"�.d�/�U3 �1b����Ep%Q��b��x��`+R*����UY��tIL p�M�q&�sK���dt�C�1(n��G�"|'���kk�-;�ns �  M�^�:!>Y�B��g7 ����^;'�zYLҲ:Gi ���CL�6"�3���T���4j��ua�À�bR{��RM)t�;�,�h�\yMD�ԅ����a�PC�2��CQ�Qql��u� �o`[�b�A$%�q�K�N0�t����8��;�:z9P����G������x"x���0�:/�~��j����
���#�V��&�<6e��vT�R`	V� ����qp�&H{3��ʰD���ݐ�(��� T<�17"���k�,-;�	�s� ��B�	��-�����Q^c�W��4�P���JW�A���7�����P�@t�ށS�z�i&�!)-6�䜻��"H� �thѢEQ�Tn���2c�C':� ���2��~��U��c�\ػA�w�k{n�nf<1��]n��j�``Aa[�lۺE����9�#� �6��C\������.���JqB��*�t/�Q(��z��j)��gE5�9J+���4U��
���:�1��� �C��u1�Z-G�_`e���k@�_� ��w�'$@0�7`8 ��-;��b����0��0�J��-��c�2�>���#�� t/j�63@����9G���;y"���9�s�r�Z����{ݻwW�b*��DyM�!Ӗ�4l���1����=6�|E�d�D6
�LhA�4���}X�k]w��LJL�<􋦛���=�\9r�l߾n��*�9��BE��>ڻ}�f퇱�C���\v�e���*�� �gq�X�lܲC��q��ߺ�z썍4*�������z%B�#�p��0��bș("�eȈ���a��6HJ�Prm68B��V�� �P|�f�8}p�t�*�yp2��*�cH�8p`I�@$Y]V�=O���/��^{�|��7*{��C�-[�T�j~~���h߾�j5���=�( ���oQ���{�2uQ��������C��Āl63��Ϧ��#�5T<G#�A�-)5�D�07�@v�ޭV�6���w��,v��U���r��^G��Q3Q�|�A����A2ۊ]�kv�y�x��x��0�c�%��g:��
$�?m��˿[+nT��_0�c������\��j�Kp��;�ݎ�B4tlqJ��^J|&��.���^�J�~���5{������"D��A{D�ؘ��榗I��Bg@��u�$�5����+k!tκ��t�zY]d�<��p.��r���jȍ�� �8�ec8ǘ�H�@{�̙3��ō�D)wyȌ%/���@�\Ï�q�X�\{���ģ���GU���#���9�x8�,4kҤ��?Mv0��� �o�4i�F��z�j��?����b����+�K��$1&��=�b�Z���ݫ�V��ѓo6�1��k��B�C�y�)��1v��]{����y!+���C�`�эNq������.sn��r���Z��v���K��������'#��` ��V�M���;)c����q�R7�zh��!e-��d �������W��At�ށ?{8��Gr������X�o� t� ο+��RE��GG���Ɵ�駺_ʴe}ҧ�� �}��a�rb}������'�.TU�~*��%������|�v��͐A��J�j5�;%�;�58��2�G�?�G[�6�d�{呻nOA�ě�E�/���U<���jժ�}P��(��D����`��r������s$/�\����儧c���U0#�Yƒ�F������J�}����j���y=�9�9 �� <�ڭ%)�$o�3H���2�@T� ~�gT�?�v��J��t��|
��)��K�	�S�s����w����ğ�#G�B8F�LI�f�ϵm�V������߲eK �k���I�Qs�(�5�SH��|Ǉ�|�\�B.����#��'�.J�^G�}�^6�|5j�tx�ii���lپC�K9��8
�8s�ףw���^��X�|{�b���0:��֭��}�`�*[Xp8��A,'�yL�^z�ѣP�(�$�����bA�"��O���f��zt�,� d���r��砥j���p#�օժ���7�IG�~��R�� �6�Cf��# B�	&��Wz�[���'��G�����P�4�㪐a>�Q�)�����We��ӛ�Xk��Ax�*Ua,S��FT����c3*x*��I(37jԨ���D8�}���}��!�cG2m�˙�,�A$aKb��]�Y O��Kr�u?��wG������C�!��`��6�c�:D:v�&�UkH�s[I~A��ٴM�1C�09������k��ɱ�1:1�R �����bw5(rz.G��u����˿�+s�l�qC5)����@P�5��+�����KW~^%G�/v���Ri�V��APJ�{�"���xY| �bSޣa��к�� tq��=�ʛ���CO�`�75G���z�!�gY=O`���s�ٿw����Xw�c�Ì'�Q:�������B�a!MF%�غu����느�P��ݐ���r�- lܸ�AY܉(Q�]N�:��Θx��0 @}%��q�3����w��˿�I�GKl�-�[��_��� o�U�=�{Q�4>K��fe�Hn�C�m@�Y5�S��'�k`E�TR���`x+�t�9��y�׃�����q�-��O�nbjT�,��1� V|��8sˈW{�ѝ��kT��$���yc�<��^�QD�fF!�h�>�vff�����4i�3�$5�BU�c��y�f�3g��"\���O�Aà[Jjc����W�Q�����b~>�.FIׄ�ﵷ��&Ѭ��>�������p���Q��vǎ�%�;�
*D �s�LY�+V|���~��H�|�ۤ(���۵[��GL�<�CbZ�(x�x��u��٫��9h���n�}�BV��N�W�@D�|q3����b��=��\�l����?�J�� ;�B�;��ўx�7[��y)m|�ͬ] }�PE�Hv���IV~�5 �y�)�x��Bt �}�*2�d��=
 :�@`_
� �ź��5�L�ܲ��>|��]���o+î�ǇW�
���:�Pm
���a�y�f�3��i����n���5w@�f�Q�PM�� �@@/�� ���@��%�s.9rD�7���]322�՚��� p�(@�5�����:uQ_ �;nK�Z�S8�ȡÐ��I�6wB}�X�?�n�im���C!�=f.�F��'�g| /�*���=%�Apd�ܹ2�����U$��'�z�7�Օ�)L��(����^\���\o�l��P���3�C"�K (=�>%_��A��#i}:IK ʰvxB"Y����/_�&}~6�us2���=���G�- "[���4*�+;�3�&��~���;� p���^����C���~�b��9鹢�D|�
h΁C�d�;�k�8?���"@0�Db���v���AD���?u§�3g.z+�k�8Hg�W����c��� �';�n���(g�aL�m<AN�Es������Qm���������2WL7��:���%��B����d�b�}rr�S��Ǐm����I��i���k��Q*$0gG"��y�KG�zշ/(�_7�[�<&$uʳ�ݗ2|��\�V^B��"��� ַoͬ�2��<���{�/ �p+1Dx�� ���Bǟ�"��IH��=�/�P��������e4��{G��~��C� y��������NZ�6�#]|�����fV���_�^y$��`��� xlr�0�DyN��)�ޘ���W��+-&��U�����ΛPMm���uZT�>��[�I��� s�+�eH�N=����jj2X���4�5�7���ډ��[7�N!���Җwp��>���q����7���3���9�B�̴@��d5@Иy���{J�j!�H�$81x����K�z6��us��I5�)ݔ?���<����S��7�P`�c�<<Wz x���D}KX����&M����Ç����'�����h�4�#k�$���BdbCK\d��_�R&�z�,���`��qz��ƍS��H9�(QA�����4��wɕ�Y4����R��r�9M���}<K^���4L6A��.(������o�<���)��S=�kM���Œ�
gHW 2w^�J�=�Z�5c�i�Z��A	��;�-���AD��%߾l�ay��t�X����"�ZO�"�A0�i	Ȱ~]�&�)EI D�fఱ���u�S?b�7�8�o��9�MO�r+ܮ'#���k5W�}T�l4����J�U�Vj�b')�x �D&\)��K��ݐ�����0�t�z�c�C�	Ώe˖�E�K��n�O�LHv�����L�uD&7h���ُ��������>0i��~������[�ȇ���M�k.w^�|���2n<�8��� ~v�7wIf��i�������U���@S	�KI@��/o!}�]�Lnh''�t�	z�K���R�㇚�9�	5n�p�#O�~K�(�@�\m�J)1O V��6{�eX߮R�lk��#?��Bē��A ����Js��v���q֟�ڊ�'R���tOj>�����S��L�г�ꪫ�J�r$���`3��*�8��+"p.�bZ�c�^p>�Ф�#�ЬY3EP��'�1]����֭�*��v"��9��X��]:d��/�G�ARY�a}(Cꬽ;?&&��N�4EF���đ�8M?���x٨��;�;Q�u�)�;��m��7����m����ތZ�l���˨Y�n���)n�ه�C���☄�f���`�̉��Fi A����9=��1 p�rDڨ���7� 2C����%�v��(�;�/�B�^@����=CL� �����uB�ނ�h��Щ��KF/���]��W��:����8����A+����8:<��R���A�	���(e�dN[��d���v�f �Z��
��U�J�;$��_P-ݣ�cҼ��H�����@�ޝ��Ȕ�㻎7A:v{NP/����E=���\�T�xX���{$���ի��}Cz᧰�f����b/Z�3W����6��~��� ����/V$������W%���-��A����:��� 2��ڧ�P� Q��پivZ�S��
�ki �������_T+���Oz�!�"�	|��ш�)*ܗ�^�i�4���f��-ީ��'R�E�F_�?�� �T�Vy����!&|n/2���/��D)7h����X��O\�F�v�9�eܻc��{��[�+��Vz�G'��e�F��0K	c>^1:�݉�G�;N�z�9)�**5�TQ����:	&���*8P�^oZ��5�ľ�X:�-+�H��4�mMl02�ϑ��>�%�ڟ
��hhG� �i�f��bt�If��R�JHx��㨗K͜(_�
��z��U%u�X϶M3��=�+�X{�l�ȇ�!%Ə�r*�j.�{�J<M��D�u�R4�T���t_����Ǡ��4W�+��]�՞��^��6ym�[$�)���O{ e� �Rf̰	�^>{��_y��Y�^Im�h�J��B���s��ݲ���2:c��[׺fu(3?���;r��'3G�+�w�*>s<V�>�0���a��/J��f4ޑa�&S:t������ʤ��Y�<A�.K����#e�΃�pF"����ԇ@A� �_��W ���T;!$A�Ȇ������͏!��# B��BR�m�*@ d�����y�A ��2|�����Ν+�֭SEL��~I6��s��P�6sH��*��k�F�٥��0t��H2ZK�h��|�@¤��Hj���R���iФ��&�H#<�c�/J�����Z ā_�ɷ_#��7YL���ۇ�����=�%�7�]y�SOq�����5�����~��{���R�GM�y���I�y��T�3T /(��_���#[�I��F�Q��Á������0  (+���!���_���N��*Ԋ�+~4�x�}Y��0I�,����v��u�2�;�k�h���ჵk������X�'��n�Z��Ǐ/�����׊�=��s��.��^��xz�LZ����Sb�	*
~VsV:�Y�72V�[J�\ N���#-\��ݣ>Y��b���5�TW��?<��n9�{��E���b� ���3��1�>[�JƌyWC���&�MMf �BԱ���A��4�f���%�{��a"��_ e�`V�h�3(�s���˜��KQ�
Pb;ԐL�_"�BL��G&CL_�X*��#��rg�����    IDATx �8ѕ��o�A���#�K���� 2+-@0�d���%�e�+���C��+?���w����N`A��q�h[�?3��>��D����f�)����a��"���Ep�G����G���B��3�J���f���k�dL[�}�w;2��uP?�<��D�H�ls��g��RFK��`l*BX���?"���Ǝ)OtDV�E�_�KP������/��W_"/=~o���*e�C�.�����0A��j�Y8�0�<����_�c�8��&%��r�7��(����];�w�|����2襮�P���F�4 ��{�����Sa-&^�߷�ݿe��a-~���>�Ah��ëCL,��?�*nڻw�2���aj#	lMN��)��o�գ��'�6�ڐ��z�Ih.J���t��.��q���\��A��3�<Sͩ(@�����v˘����ɟ��%JcH(=vX)����x��$��>t��^��YB)�PRU�vhD��CƎ-�;twt���YM �O��P�Z� ����K������%���BJe1&D��7���`���f����/
�,6������.{��P� Oi�A�;@e�}��[�  G�<۫'<��}��u�u ���=�"�G��r9y�ϫoJ��ń���M" m@����jY	�
 @RgL�:�W|�]w�0�W���W��aÆ)�M��H&2^L%NVIG
�ip�z�5����됒���ŹU�_Im�YL�SyN��sW>0d����è�#S5^!{�{�x_,^�m�ԆNl1���AOh"#?7��ȃ������x���ȕ<V���,X�\ C_��Q����kY|��l�����$X ���6��Q�*��`�Yp52%�[��w�w�tܺ��乑Rk�� �C	+�	!������@��3��Q�K��ەR%^�2TmT�^x9��%Rԃ��J�^}����ՠIuP�V�m^�aj����}�fL�>�֫��Z���n��{H/�w�Qa�O�"�a%�9���=�,��=J��x��J�a)�+J�����(Q��|ڒ�W�1��l��q($��G�d3]�.r�:?"��x�&1(sp���ob�����@�}��2t����C%s(;H�z �*"@0�oǏF�g�����U%ේ͆����du�\w����3DXMVS�` ���d��c�iH�8�cK�UuǾ#�F'8$�B8�Pq^��8)������	�o��J�����Ǆ����~5[��ɺ	�� e1g�W2��E8^(���Ży�܌JX���CK�\�^��(�@-]̤�����k]���+��^N��_:�Ug2 8��d�3
h�x)c>_π1���B�:�J�9$�lB'6+���^��B!l`���r�m��!�m�"�����p��g�u L@�/X�ld�Od5ţ��-��X�n{_q�D{�(`�����b��d0XM��0�X��G@�3��\��h�J�6o>BB^)򀄆<%�=0�n���5�z�ld��1��q�%�
ޤ8WЫ����+@��vI6��o���-7�FK�H������T ����	r�;�W\!)))*|�y��ӦM+�Y��p�>x��� *��]�.��CK��	�3f�I����r�<��3�zd��ySbU
�|�\�c%D@��GF[�`����V���d�Gu)v�����dń]�Lu���=?$<�&�oCq�\�r�����_-g4n �hV�s|�Q��7�X� 2��.�F�|�J~9���d)r�!��+��@Z���}Y�Jj�˩�!������	��j�h�N��O��aFU_��E�7���x)t���/ʄ�B�k�n^5eH��y�:�g.jٲ� 0~�FT�:�]9��Z����Y��_��9z�
|�xc
,��ر���\��5����J��Ӕ_<�2��IR���J12�T�
������	�k
���l�#K)���ħ�U��58hr�P�C��@������E�d�fBP6�ۃ�&x(�kՐjժ*c�l%�:�+NԒ�k�|�Y(v��`��:������k�W�P�L����Q��3c��$*��X��u@�"Pā�(.��Йn�����D���� q޼-[珬T$5H�S�L�F�N%M�i.���N�1�M���:/^�F�7Q�s:z�y�wʹյkW%��97r�H��g��S �s85@x!��v7�9)�!E�p`&��"�������� 2�O�ʒ!(a�5���@ <#�!����/% �Q+~���
ކ���{=A�0�:ߚ-P=0�Fx��g�������p<7�=y+&���c��L	�e�� Q� N< �PS׆�ǐ���.��o�ԏ�W�B9d(e̞=��~���U�4AQKh��G�(꘱��0Sd^|y���+��zL��~��G�n���~'d1E�<�5c��'�3�}�!=���3��7��X;@FW绛VB;j�q�B�D<V�NGV�l6
/qS��9 ��^�L0�.�ؐ5T�l��0� V^�1�UIZ��ը��cQ 
��yL䳪�ǘ�B(�L�����@ƚ�b�gA[Q��� ���*�)(a1���Z`�^Aąv����e�H�X���L���K˗/̪hn#F�(�aN�c��}�u��.�R��$�Dy>���Zˋ���S�\`rqBQ�Ҵ�� �����Ц}���!��'@�uk>��īv:�t��c�����@H��
���,Ey�!����8TV���t���9A~Gq�"�}X���.k��X��+�a'��������AС����Y�h%nBC^ĉ�8;�f^��,?[�z�w!��
��FF�)T_�0@�{��{�����7'�����Ϻ�����Y��)�q:��F��{K�,y��%�����t�����kM,��Z�!��=J��x�|��}ɬY�J��HR3Ĥ��H"
�<R�/�:�q���骡< b�!��P���� $zc0�d^p���=Ve�m�ͦ4V��n/>o�*��[)C���?�<Ȣ7��,  �<���y�����)7<�X��2O�+`�<	O�o���G@�P�#�M^��'��D�a1�2�a��k��\7{ؙ�<T����-Zԁ:��:䕩�e��+W
@DIj0\��\O�ED���|6����'$I͂��*�� Q�S$uƗS&/���J����y\����A��El���������wa�o����X�H�:@H�$�`�<�֝�b�%d���N�=�H0�Hh�C�Qxo1ՃP����o��<��!��]+���SW� fQ� �f��1��༮�P��c����;�Ѷh�W#}�� j[�h9�Q�Z�Bʻ߂�޹s'��~lI�i�cj01���0i�a��H�Ae�E��8��B��K|�8��ra���.�w��Z�FCL�9�Rg|�X|@X���T�A��2̐�p���� ����6q�M�o_�G0��{��?@����U$U�&����`�ȋ�&��*��% �܇���̓0LD� WA��
L���x'Sl�3�gz0�i����w(.v��`>GP�5)����麘��� PIͷ# b �L4��j.�c ������GBs�P���
HyO��ѰRY����<���������2d�ʤ;��I]�C���O��p�^�^T2���%!�P�R��'�<�ȱ0_��u �/�� 0�0�\-�@-��S���\�ab��(�F�	� /<����H��j#��Q�����"����W/��.�*����J�o��,��5Ө��P+��,I��!�E�¬8K\�IF���=Y?�����Ax�m��Q&m�j.���á���|3It��sl�ʖ�|�9�Q����j�*�y�����zq����\�(@��4 @�N\8�%V�	CO� Y�:�H��߱�WH{��\p^U���Iӳ�����NU���E�>7R~�u@��i�ϨWK�gvU!�B��+�%9�&={="�p^:G��v5�lؑ��q�e�����%�~�^�t~�EY8w����X��Sr��d���T���2h�B�|�ʃ0�k�5c�M�&[7��3�H�nC$-�%AjY��^�>u�I��'����Pr.�!�2�dIm���8gX����}n��N�8��zi$qJ)l��x뭷J8��B8�`GE4N�U��q^Qo���N8��,�c��IH�(@��T�Jm0dҵ��SW�;�<Ų��e���M�{�(3�-�i��H�;�Go-���y(���V�eԛ����M7�"]�zT����L)�������Kn{V� (?��$Ha��?P�"_,]$��89^�%藛���[�7��e_L�n�G)��2�i���U54������8�
d߮����(oe�g����ó����ɂE�ɸ�S�Tk:H�+�|3�A��]�g�=�~VF����}n��ѓ������	{�tj�~x#�k������y<�-�d�=Sr1�=]g��\�D9��O`�dN[rKڴE�2�s/����^8�ַ\}�������y�>x@z�f��g���v�\z�����r���a��W�}�� �'�֛���o)�i}|�uwK-J,�"ϼ6U�_�YU6_м����t�c2�㉨c����d��%/; ���rC�Ge�S������z����=�姟~�X�������e�w�d7zkw~���;E������^�p�<��8�͑L(,�t�D7A��S�R�R	 Q���3��Ij���(�!;����w��~؋y�,Rҕ�:��j�*A��6�bj�����:��#N�U��1t��@���ښ[o�Uu*��
2�a����9q( 3 kD0�Y�`�Q?�J���<��Qy���ҷ��]PC��G�,���f����;�Q�jd0�}���sd���rV��m#w���4�i���f���\3�5��uw�A7	�
?�U�.#ޞ,�Y2,�9����d����/���7�5�>"�-�*�_%q �_~�a��u��
��Hz�\<VQ�G{�Ȍa2o��2a�L��=q�X�5�3�3�#%]��� ��AI�ʉ(M*��y��5 �g�����l0�UA��.� 5�^| ٓZw�� @��}��^�ڵ��l�H����(@�Ґ�#v���|޵lKd�C��L���K�LY�0 `X	�����vE�b �ap�˪�ߕ����6�ޓ��ޑ���`XE爼��p���X���F�j��#^Tz9�K�yC�֬/o��A��~(�V�@mD�!:���.�T�<����g�������bx/�Ȱ!/ʵ�=.K>� E8@��lX�Q��U�â"��H�&mrg�G�]"o��,2�D|�U�����)���/��/����>vt�chYR,�cUw��uup%��|(���!��)_Bi �<ǁ$5�ΩFA=z���z(T��N�h��)I�?��4UB	HT�,u�(����V�D�
a���3�x'u�B�+hj#�:�hE��N���,Dfdpf＜�R-1����8�J������:�d/1�� ���^P�i�8��R51	}'���U:��A�[��W�0qV���edA���� ���<��/.,?T�G��j�V� ���e���	i�fVb�X���D
n=�'�s��U!)��!S�`a?x�,~�jN�jpڗX+�2yРAC'O����<� m6r��;v�{ｷ$��܂
���.��'C���.P%Xho��ST�H ���  ^:ea<��y,JdP�Ԋ�:-�j,I�cR�p�1�`e��4� &��A�R���k�/Pշ(�� \�0���ҙy��P��1�CX)��4D��OM/��쨡H`�Z����=���ƕ���������l(�cͅ�ҋ"�TI�@!i��i�в<��)��*1�gU��	Xe�\ُFI��m�~�<�"�$���rN�����M�Ӄ ��٨Q#�~-b��QNS9zڿ��3G��oZ"Q��j�>��k��hy�/)��F���-x�,~c{I�/�Я��9 C^�+�KVר�Ǹ>�f1�on4������6��7�#^ GTT�L��?tX��o��`o nly����) �PE6��"7z*X��b6����"?�]���>�����5��Q˕����,[�d��xfx7,�c�,�@�N�*"+�A\���{�*̓ ���믿VCǇIRs�z�1/����%6/u��A�*�u����64)�k?�̔�)+�9N�ޣf,@,jA���XlF�ji�;WF��%��WS��=*^h��x
3`�^�C�U�(BS�曞}�:�U�k���6~�q%�n�ٽ{��(��U�zu�V�����T"N <�F�g����y�V��ʍF�F�E��+[��F�E����=���o�.[�l	i@�"}�!����H�ƍ dV��,�-.�T���,?�9���%�7U�e��4Av�
[%���&@���ۡ�T�Žա����(pT�罢\�JDPp!B���7N5:I��M�6���M "f	��nCg,{#mʢ+� �����c��)�9l�)�˔f����e����+BW�p'�C�/,��~�~6�A|�ȑ#�D���!n��;�����%!!;*�U9`�	$v����!�)��N(1=+�qpb�{'C\!i���J������$<�{��6��+H@C
���~_�5?[�{��x$'�^>��� ��J�� ���{J������'�1���&=�"� *�QQ�ož����.�cØ���0�~@4+�o����bj7l���R�~~;�\ى��0O�a���2r`?�w�FҵSW������- iMI����U�ғ�||�;�q����T=9�f� ����]C��q3@��>��(�g�����7 ���S
��Y�zܺ@��@����2!� *u>&6;���dD���a�C��(�;y�$ծ#O>;D~�}�Lhe����4�P�	 �ā��A�������4�A U���(� ��!����{�X�^���<Rj��I��v �DI9
' ��������Em���>�~�!HАZQ �˕���#��S[�w�"���R���r�3��4�+��X-	�P�:\�U{�.��\e��J�(��  F�I���H2H.���2P$2 ���	�.�D����E�P���S�Uu�S�-�0��ǡ�kaQ��;I�7�#m��ʺ�� ��� �Q
 V�J�I}AeT���?�TV�R��+8�z�B�W^y%T���(.-�Vm=��Z7�_&L{��cx}�����g_����ͦ"K��D��S��g0�Ԇj��D<�,��C$`Ǻu��*���_���5u��WR�-m�0�R��
�B�@��8Η-�g  ή)=ǏV��7>�n���0�|�5X0���A� #�`�)�3j+��GM*�r����Q]�`�}�#<RO)�
kµ��>Ro�P �N�.��U��&����lJ������6"5�J�)����<5�iФ�<�x'�](W��q'H��AR?W���>GJJJ:��zq�Y(G=]��U��(��_�>�C���q��g~@��ZH��E������T����J�W�sC=����=W�"@��դ5�0�=�ܒ���#w�u��~޸q�٧z�g���5@��ˮ�~�/m�҇�����P�^%2�3���q��եG�n�u�2���$�� �j�=�4ֺ���d��7`- �����
�7ۆ�I�p�;@+�+p� �
WN� P`緂�<���� �.vJG)\�O��ނ2��T�И!2��A�r#�|� 1r�D�۴�<��Y}0G� �����G�͊0T�O����,I�.���g�U�� |����Y9�B    IDAT��p�5�իW�P%ރ�E�6 ���R��[dKI�o$PDA�bϚ��9~����32<����ʐu�޽墋.R	'�?#�^{�~��#��yYܙ(@� ��˱���4mi;�!�:R�c bz� �9�b���X�5	m۶U����H�5޺us(\Ģ5Y�Dn�� F����=w���E��g�d$/�,��߇�������6�����_"�w절��Q�Ϙ��n6�Q+z!`"w�W���ݯV�{v�,�S�H�8@���� g��ߒ手d}X��i�ʚ��l���
jD���b����� �qb�!�By:Q{:�D�_�����s��1f}�*-mE�{��L�݁{��6fzNh�Y�'5X腆>��Q���@{�����n�ZM��A�[�2
��{�rq�E/�M[�X�)	rK�Z��;�� ��b�����
�}l���'A�.]�U�Vʸ̞9����D�**b](eP�ΐ�x�~�6�S���e����
 �@.�F �� �Q�}�ͷJ�֭�qcǾ��AO�P�8�p��%@<�DG�϶�[d�дp��`�/1n��i�4�A��Ɏl�IM� � b�4�Ɂ&1���o�:4��{��#@0�T�V��p�&�y/4y�5�� ���+��Y�В���0SşR'��"�4���J�'���k�.�֮]+/���ynA��EYܝ(@� ���_����S�.{���^��*T�CL� � @���Eګ����8x��-[*�x��I��?(�j4C#Kg ������h?z�ȭ�oUW��Ӆ2����*�<�U�*�΄�o���r>��������d�����,2�"�TD���)���;�"{S��<�O�ԣ�N�z��~��  BL�d"@(�@(k[<�av�]��3�q��~C�(cʔ)��0&����8��]���7�L��D�=��ݜHcnҞ����V�/�[�̑�B=������CO	ץ�?���i��,���& ��eqk� �k��7^�N�pѳi�?^h��� .GS�NOI��C�(3���S�N(ZL�ǎ�U�}��M��$��K�b5��4����_{����_�����Em*�� ��������U�w߮�)Ӧ*c��#�Yߡ�h�������G�*Na���28m���02�.��(���M���01��D���
 ���dA6���J�80a�ѽ�Q��[n)�ɡ7�p!�~����Gz��?��A �p��y������F*����_��Ӊ_42;�s�㫲1ޜG�zܹ�Jq���>s��Qi����w��6l޼�����Q��5@\��[Ӧ/�9u�ㅆ�X0�J8�p����bj^[z�ݣ��W��aM�E:u鬪�9�N�&��y����g�5_�(���*BL���ۍ��UyK/�s��ƟEq�qt:�$�YP����&w�w�"���nU(f��JcU�s�=�g�L(�����c�0�s���QAd?��( D���@��O:��`�$h)�>/=�ց-���7��AdB��{䪏ફ�R�ڸqc�S�� ��h �%�J�*�:���o����Պ��aq���������϶�'�"��S^����^`(�H �#x=zT�͛' �K�by �zl�U��_s���pi�S>i_l�š�����������7�M�W�ҫKwف8~r�*�jg����x��Sr�a��üfggD�(�K�x^�*�c��6��57ܠ���-[&}��ؘ���
'zO�a�MvHw��� a���+��m��t;�2m���+�-T�D�ˌ�� j'W]~�<��QH��
1>B����Mrss���;a��9��<��m�t ���X`bn>@� Q�j�-�S�UA�\�� �Sw~�pG����"IG~�F��ScI.(h8XKѠA���x�5DrX�>5萃W��oj���?��^��oM��rס@�J�o�^���y�Q�#��c;vL~��%wC5.,:$۶m+�CQ:.2�I�J��!�����F�� Q/�O��ّ�>z��'81Mb2@�4�c�q�42M.:+I�͚/9�R��+��&Y�h��k��O˅^�z�L�2��TO���;Oj׬..����r�����F@���]�d)xa�/^,�?�L�@��� �x���������ȡ��H�o�����9�L�"�IUC�*�T[-je�k;p� *��r�5W����-1�v:|��4Db��zv�fҨAC8F�����J�Xy��Y����M(�	��6d=U���2gH��?��������&�#3Q�����o;�k{��wA�C�Åuz��ٳG�����)�ea���О��2䢎+y��Z���k�͍���#�(����BO�c�駟���]�v�������]E�C�:���s.Df��1¾k��tIY�Y�z�O��a�P>1Ь�ύ�4��+hOr��M�*���0�6_��I(�7�ʈj	B��\yoݴM���V�j\_���@?i٪��\����#��J"��+�ݻ�VɱV%�g��ȱ�\��Z��g�H:��N>_O���;d���v�d���rJV^�B
�_W\��eym�.`�8 ��m�v����$��S���}�K^0F��Gv?����,~:>�!k~ރfI ��bdGl ��6�l�3�R͟� B0��\n:n��`O-i�ЅO|����M#A�N�k���X�I��P�V��T��?}�g����$q�Mc�"�a��J`x�'J��=ԞƁ�Q8V�Ü�Q}VT�{(^�)�O��c�Z�_{W%Uu�_-]��� �(�@�F�H$��dU�d\2n�h���G�F�D��8`2NNB��pK�T�5q��A�Q��z漢�{]�g��X�v���s�tu�{��������5�1��\�d�Įs���T����@՟��[;k�Mˎḩ�����}�
�6�@
�6gf�ӈ!aU�V���"�d�7g�d��`�>��Q�xSck�������pmѷ)x)LP���B ���FG ��X�1x��w�+ĭ.#�ah�Ӹ�,� �F�꛱��B0a�(DC�Q�tm���?��Q9��1G����<��)�DT/��cF��B��Cm�5��1(Fa��EL,F�j��,�+Xri�W��v#�Ң�o[���yu�������6D�>��Q���)����m���i���I�B�
��~�����]kE};����>���6w�ڽ��&M�,Z��S�8̩5��L��N�܈.x�՝�����n��)X�M�9�c��bF�"�vuDe�gƚ��6���j��$���S�2� ��y�J��W�R�ZF>C�"J���(��U%j����y��&��K��<�j<� �SAQ��-�*JyR�7!{j�忏>"��A_�*�%X��#��Kn���(��&p.��ы�ŅfO��u�w�[h
�\�bp-Rdd���P���L�-s+3��yn�98x�>��}l�F��W�|'8s�σDYe�����:*`���3����RA=���I�DAQH���%Ek_����]LRWm��F��c>
�b���X�&[=�+cԆ����[n,��y�3g��W�kA����c�>��v	�Cߏ��)�Fˮʿ&��3�gl?����&�%S�3_�玃���v�t`ꫂGҧn��y;qQ��<x�cfߣ#�����箾���������\&�OV�54�'�0�B�6@�2:�$ �uDn$z)�͕6|\1n0y�]C��7w�>�<RtC��\F�H�WI�4�pV����`�qG�ΠZ�9x��U�^4��uY� ��(w+�,ߠ�!!��4������;�k��(y����/���w*U��Sy0O�+Y�E�!8x���������ڪ����]4%Q{4�ҤL�QR�_��G��\���BS4�8��jm��mx������$u�FgM��?�O��j�(��g3<��ڂdp�E{�G�jK� >��ओNj�����?���R�[f>37�-z����O��rWAՓ�$�w�$�B��7[��љ�)|>)u��K�)�NG��������'��_�At�Oo~��_���3���v�l�,�*o�TqiIkssp#�F+JK'��EE麦��lK�bxY"(C*��wz���q�M��S���:��56�:X�s���kH�c���N�Z��{}|b|s���Dy��X�Nc����<V��ה��)���ϯ4��������+��q����lK�,��j�	��Bo���A=�-�!�O˟~쑱4v@/��~�ÅK��x���ZQ
��$Y�ZB��u�9Ըc�Qy���l"�mMBM��,+Z���_�$aX?�� Lp�n�����1�:���(�BO5


��2����&Kb��g<�^PQ�5kք^ez�-���P�S�[�.�\f�ɀ�0��n��`�����[om�U�;�q{&�����7�pc{g�����t<�ct}�g��دo�i�����<���+��ۛbE-��!ٺ�\,�J' ���Xֈ\	�0�a.I&�Q�4F"XSɺ��?��5{�:q�,<���M�cϬ�OÊp,��ݛ���M曇d[��~��o�'����A���s`&�liNA�W���<LZX��rH�����!�g�z�qGތ����}v�����[ْ����8�ɖB��/��̃#���g����;�N<��,�\��[�:}��9����`�nB���V��͉xQ�7ښ���\6�L�q�|K�8��)M�����B�ɋ����:7|0
*&>�e�	��~dT�1""|�m����G=X�ืij��e+F�Ì����/B��2=��$��ۈ�(�)�I�k��5�ѩ��fS��F�T1��;As���Yj�μ�GÔݳf�
�`D@�W��?����O����>� �Ĵ_��u���n��jk}��-�쐡U#����B�t/6/a�P�B��i��t`�����-W���`�~����J����a�h�����Ft�/E{�g֯��[�t:SY����xM�_��bπ�A�F��C	����MH�r��d�ǕUeO���CR��8Xb�dXY0��muh>򖒙n�GuT�6cb�_�v�J��w�}w�6,�T�7�F+u�Yg����}�߈�|򭭶�-a�T�nfK�W����:�@�J�cw�uׅ��g�F
xfMX�zuH�W��N�UT<����E�۵����ǚs宻�jwV Q�:\`p��sV�H-��m㡥Uj�L�vH&S�E�?��rh����%(i���ޣ%�[Tp*5��2*ؘI�e2�٢\��bhc��d���N�`4
�4&�.�6Ta��$�C������-���ѹ�������4�f�FԔri����u��EL̿�����/v?��g�o����sx�]z�a��ET+������ێ�H�j'�o��(�����.�D2�k0�&+6c+]�g�!{�f1���	�y4��τ�^{�\v�e��lg�t����nhSb&����{�n�;��/�<T3Z9Q
|��H
��s��ɜx}�����_��T�l�=��j��n����MM{l�m�'�o�}EY��$�>tT�����a���Rגn�n ]^�IEE�UL�.��8'��5n�ڍ�c�t<��7A`��9�yt��9�Q<�?6���"�;cʐ!U#�����Ї��q�-��3�U�A�M�Ɂzh�H��QE5�!Np\x����S�PpPM��	�#1x��1��]�yPY��	��?Ӄ��7o�l���(�`�^I���Q5de6I/%�
��|ZF�C�ј2eJX��^Oc��a�*�/�y��.�k㮃���WH$\T��]�\g��U�����ޫӥb�L����U�A����+ә�T�	�gY7�;Q_S?���al"��!����S�w���d��iܺ�9�(����lyI9Ie}��d/ihȌ�TW�aj�d<5��j�K8�Ϳ��wULps���*�E��m���	x��^�@��z%�M�?��� ��@ ����k�Is7��}�ܹ�AWfs����?�A�B�\��q����߮��H�o�ޑ���#��MR �*)�Èx�)Pؿ���X��S����vT������}�{p��0תa�h����ys"��ݑ�Z,T�T��k!��A�v����P�'�\z"Vi��c�5�_����_���������?{8uG�����J��L�+����A;�!�s�k�6nL���D,Y6d��pν}�W�5;���5�S?�S���c�@�VywB�p�&1����9dԨQ�Ã~�n9z��` �a((8��g��{	W��1E�U,#r�PnF��.^=�:k^IW�]�|X$�8f$y~oAlXH��huI���=��vo��Z*�[�1/�Q/�SU����7Ǝ{>��^��-ȵ%�2��m�	��DhmQW�N���1��b����4TW�?�bl?���7w��Q<h��[�V� ����СU+q'a�/�sxSS펛j2�/K%E#G�ܛ�������O~�ka��ki5�`.Y�$�~�p��ϒ_C%xV�otu���3*�ðK8����r�a��G�Zz�m��� Ha�=�n�$#��w�0���`d`.��fD�p�����fD�I
�����ڂ�s�;?�C��c�e��}��
���X4v���5��Q���TC��hˠ�{����6~iY�w��v}�2b\�v��'�=��|���0�� ��0��aBu�B�*&,0��q]�⥥��CKJ��y]A�9�jZZ&���O�r�E�T�a���94��_Vr�Vo�g�#��
2�0��.��@��PO��$N�0��3	�"g�zx��ۋĘ0Z�xq��0c%��Z w�O}���#@�9�$
�����t�*F#;��������rk�}��Σ�>��ӌ�Cп����Ǐ��1���*�Ĺ���D�����bb9v�A��@��������1���$WC���S����j̦�=��c�H�4u���dQ�5K�5��H>�������Vݘ�Z[W�C<V�,�l7���8�.��������<��`Μ9!.�Z�jn9��~8aL|	w���ܯ���f|�ʓ1�����d�_�R�P��˒�ɋi�L�0�Z�{��C̩.2�4�rQ�o.��;�1ޅ�b������XQ2J�H�}�J����H���nFZ\,pWBu��H��9����k|q��%�������B7Y�mi9��m�gL�*���7n\&|�$��J��TS8g6Ҙ�յ;Ã~��U:d��z·����x-���5��xa��.)4�J��
WW����*�{��<�*s�����	�`����ԩSC+$�]�y��2�����ɖe�T�ֲ�Dw0�ѱ_��4$[փ�=k�}��,��j�SAԓ,��ci�6��B����7z{7�7����>	�H��w�_��z�@=&	�����?w���W�!FaR��j���e�g\<&��0��M�0)��T�U;8�k �
W'�a����K{��g�w� `s�k�S�s')P�S �˰ʿ��������꧰a��=�~��N�,� ���)��2�㇂��� �ٗ/�-����W�]#(�	3�I!�'�a0�т�����V9]\-k�/��$#��n���T�k�+��N������Ci��J��[ �qX��8L��c=������J����� �p���]�4�������a�k���w1�R �)BC�ֻ0�]2P1tݯ�¢����� 0[ �����X�
���J����L�f�S_�� ��ʂT/1�_<�}!�0�.��۾l�qfX7Ae�x��5u�]�H���5ym��l�9$z7��{5b���믿�^�!L��+
� ,B��aެ���$`ӥ�#  IDATz�~!R��x6���s�s�����V�:�"�7w0���ON�@����+��w��{bb�X�	V��u�ߍ�?����X�zL�'�W(��tY��}�(��k�)�9���n����F#���D�wS%�/��Y�
z����[�r<��������V�&t)���_+&D�k��Çy��޻�p����g�٧h*l��X� KU1��%9�m�*@N��c4U�;;�����Xr!�׷�����#��@6� �9�w��~�\E�s c�W���F��1�]�A`b�@pBa�4v�C{���W��H��?V�;�s���޾���ya���/���l�F�V��$< ��}�b!���a6��ܳ���	q��ɓ'��m����.�Φ��J����K�����S�X\�m�2&�)d:�Pm���/�>Zm�c��(!�z)�v�-V�8އݯ��O:�y��89N\X�٠@�z����#����#��ys8�~�#�<@J�犕+W� z�@<.p���j��0���?v�OL�*��>L�]
A_���'��R��Q��� ��s���B5��ԓ	휅I[�v��C]��*삁�_��x!j�l�M��@��O?�=/?� ����詏X$L鯠���k�@X0{+�Q��e��g�WL����z)�����K'a����������*��f�����?��pc��-�FN�ChS9�1�R�	%1*9Ӻ�Cd6#ɩb2B��s�[�!��F)��a�XLr���3~��G׃����|�]��a�Ξ��5
nFh ��q��q_��u��*2�8�/k0�#aFӖ��� ��{�>����sRΐåF�����w�E��r�̸=Q�\2���Z��6\bTs��E�)���Vt��.���3�֨f�<��E��p��/��ZL�p:MC۫���?�U{51J����X�y[bK��V�j�� �0�x?ΚJ�Ls��cPԖ�@�1�z14��^	^��Дq�p�!�t^_��qJ�)���.fr�M�j.Ʒ�EN���Bq̓���n��B�2O������D��"�
V5~sm�Pa�ωYh���^�r��	rl+4	�t�-+6ѐ���B�vN���+�R?2t�U�����������6�k;����,f�9����
Ƶ�p6�^�^������)5�a�����(B���CWz0���Eǈ3E+�P��gL�N��k���G8�{֯��~T[!yXf��)��E�kM{�[����]�R���m�J�P��OCZc׿��tw�m�|���+*�Wݞ����­w�����ַ�:Q%]��I���Ͼ���O���և�`��,��cJ2J����^>�A�,@�֔sӒfu�u}�#�A�\��Z֯_�ݛs���F�]1
1�kwu����I/�����AŐS���N�U���H�i����iҸ�m�}(��5��� ��i�U���1o�VnXL�E_ԝ�~��l39C�PR��)׀.���;����.R�����rR�����j�ͩ�8r�UN5 &>���^�+M�^G�K�
G,�<y#5�[�p����M��@-{C�����#-�i7�+��*֡����[�1�h�Ե��L��Ǩ���=��#	Ɍ��A]=l����JS!�@�n���c<H�O������N�]j�k-c�8k��{����\��s3��Cf�_�f���d�/z
����_|�n]�=1I.�f_[�D�-����:*(��\�x��G����bm8N���w�@���k��7�v�:R8t>o!�.�Ev�Sq�݌L��2���-j!���Z����F��E��o2�c㱃{D6I#U[�#���x����nG����ZUF�,ċ�=��}y?K�Oz=.O�G��<abn�75�!���֘)�C�3�i����#��t&?�
�tF�}o�tY���Ŏ�<�����Z��_FOK9"S"�Ȝ����IPaT��'�C�e����/y��(l:��7����Jj�"=;�3�{�D:0LeY��F�]�������<��V��u��g�k�H�S��F��r�:�����R��_w@_�NZ��V����\b����3!Պt�:hv.��ڟQ4K�j�=�0�t*��	��;h9pVc奋}�m��܋+��Kۍ���!�n8�m7�54g��SE_�T%pC5	@���b�����8?ݎ(�Žt���>�?����X3h��)z{�:d.�7�ʹ\�
5Y��!l��%,���?�d6~]�j������.qzyP4c4j�A&.Dڤ��,��Bp����2U�;@|�1}ﶢ ��ͱ�sN��&��*���v�w��En�X\T^@Or���a���_=H���ll1����Ay4�X�=����t8�mke���cC�_�����bR�h��,�>�bK�'��Ƭ�0~(D�$����<�q���x0�k�
�h?d�6�傗�i�U���)x+��a���,��M��AD?�>�1��m���ff��Gˣy�52ŗ��?&�؞KI=��*NhW�����F�����]�XM]J"RV���SL#T!�O�wL��h^̭$y��جY�������nX��s�CF���W����Þ�	ǎ�t�(;�h�K��aӽv���|-��*9����x��
�`�J�z|���!	ą�� ̲}�'�`S��}5Q�4�"��d�X?1����㖁�t�MTó!��%���sӌ��Wk��I�7ș2V�VB�k�ַ�g�i$9���K�]P)���K���Z�c� �����҈d�j�P i�y+�e)���&�>������5q�`J�b��Z�(S����ƍ��%|ΣI��罒8���q"�Ͼћ`N���t�Nl���XW�����.#��id�C��]4|�o�ޖu��w��ޝh�0�p��M3l���9���#�E��������+���M? �I5���V�H>Е�(��[�V�AY��+3T���p%ư�J��:��?���	��ve��fOZ|��6��6�"}@7���$�����(E�?���D����Y��2��8�u�����3��|T]sq�,�#{�E='����o�W��T�N2՗���ea�A5�/��x��4B��E[��c6�7��~�1���a�u{w[�Ak�렎6�s:�:*� �Z�$�Ip�58��-c
�J��W��r�8��z�+`��@�����o�#�X3�4[+`V��� mt���.^��d��.`�q `7E6w ���Dl�ѣQ#:I�l~;5A�N�=nϯ�&��N�K��"���-U��U7�3�Ϭ?����?�վ#2jwGG籐�?�`Se�M�PK   ;7>Z1�o�b  1     jsons/user_defined.json��Mo�0��ʊ�byl�ܪ�C���*��`K���*����M�@eJ�NQ�~4̾c����e�л�[�j߸*�f?]���	7(�~؝������������O��on[�]�	KK{t���.,;����z��*l(�-k�+.�ֹյ��n�e�m�	�SM�[/���^��t}����ı��LēC�=�;�檩���>k��K����m������B��{�_��4\3��xj���C(���>;��{�m�O����pE*N[I)1PP���MS޴]����{�s���v�[��]�}�g\��ܼ~����O��廐��p�k�;�Ǥ�W�͙�8��w�;~��jػM"�)olӄR�n�6��˲2����*]��i�6TՈ���S�Ή�J�ټ���̻*�%���!�
�b�G8����O�K�#���9G��"ݛbO��?W��d��~�������.EѪ�Eɔ�MiU.��hU�;n*Kei�2��)�E�Th>�(DH���<w$	 `�)�Oi�(M�M�#�Ҋ������O�F�q�U�o��д)�5в* ���w.�꼆���;!v����2�9)����he�g�Hb�l˔$����j� ���_��g|B/�g|B����)4�+,=B����=(�īE<`�׋xt(�"^`�0��ȗ��â����Ei�MX���(.t�e�_������2|�c}'x4=�w�l�Y�����8�X����ֲ�C�Awf��%3]��'�zo4;�𭏅���}��4~IX@˗���/)�?���YFǳ=��iG<z�k����X�',>�Ԋ͉���ӛs�x�����oPK
   ;7>Z[��=  4�                   cirkitFile.jsonPK
   ��*Z�i�B�� �� /             j  images/8f10cd51-b334-43ee-ae1f-f1b63d43b44b.pngPK
   ��8Z�=�:��  � /             t� images/a3896090-6cd9-4aa0-adce-88a16a68907f.pngPK
   �8Zj˳���  )�  /             M� images/c68186f3-7e1e-40af-a8fa-ebb36c358ae9.pngPK
   '�8Z�ڟ.�M �R /             1s images/dcf4c277-9ca7-4718-9875-b39da06c9102.pngPK
   ;7>Z1�o�b  1               :� jsons/user_defined.jsonPK      �  ��   