PK   vm6Z&�@7  ��     cirkitFile.json�]K��8�+��I����� �����!�0dK�6Ʊ{e9�� �}I�ݖ%�.��~`���G�b}���ҷQ�})��٪*&_�j=_-G7B_��*���K����|9�W�_���~t���׿?�����jY,�IUR̴g&��8��qZL�؊Y�j��*��ht�������.��
���C�g��dF�c;-�q<U��uce��gqe���x48�LGE��xlK�c'�,���,R3!
m�8q�6ܗ40�W�����ri`�"����1�\g�u��r�)2�FF��[@chl	�	���!��T^�nq�qa��)�����"�!���v��8v��ؔ�O�%����c)�X��4��4Z$h�Ȑ�2M�J��,U4�e��*f�ljt��Y���r2d���d�4���dhH�ɐ'�/2��ICCz\��
ih�+�����DCuxd�m��g��2\���B4���C������D�9l(����$R���D����~��A���W c�46կ@��l�_�������k	5��l!ڕ��2t�D��k�2d��Jd营B�+��CʓhW"C�tѮ�V!1N�+��CR��*C.~�)#j� ;02���J��b@X#��K�j�<���%- ���a���c��j����p�?E�����d��X�ĞJY�T4�\�����R�e:����,��"��vL�i��i�k���!#��I�L!d���f�E��<������Iy�^�♴��D�lQ�Yi��)y����r�bE&A�4(N'�
���E<��A&[AQ�H"dv(֥J2�SE*C��N����%!tJs!������>nPC�T�)�K3��>����Y�����@-�����=nՐ#�ǭr0��UC���j�!N��tڪ���+'j�n���&jl�f���+&j��^�ώ�%j�V���N���:������"5jtB��8'651��dF�$�:�4@�,6u�-� 	NE�PQ,Tb*���a���P�,TR�1������������ÂĂŒŒI�X�X�X�X�X�X�X�X�X�D19@�S���E��TNn'r��rr3�$8��[� a@xy�{ڪ�H�� ��UC��TN� ����9@�S���I)C��B��TN� 9�����iIE�<R�~�.���#�y���F����yU�'�lV��r����|�2,�qweX"B�@�
�E+l�@h�|fʰD)2�B!���D�9���	422�
�J���M#C�jC���}:$��P�K�� ��/"��zLe� �����@��DNC�5
9o�]����h�7r�	��!##�TخFF��4�ڎ�w��PU|^}q�P�̇�On�����ѱ�N�@_�a���0�sb��@�3@���3xw��^«�' :W�y�>����� �EC���W��_w�)���O � �	�� .�a�a
�[�0�;d��$2� ��M5��@�"�@� ��ם �,@�J�WfU��/�R��~����?�����h���WF�K����'���r�V��!g�xw	���n'�f���r�	�O�M�O��͚���@���ܡ���M��5J �@�d0CRT�:5<�b�h5*�%*�倐��h@JC+n�� �8��C������/�#DN���9��; 
�Irt�\@����;䐣�}%��1�g=�u����\��>�~�9�H�#ʇ�'��?Â��Jw�!��=y�C���>�өiۅ�W�!�<<�\�!�Ʌ�&��6�5ɹ�r�C��"OTL����z�I��&���!zJ���9O~�y@���,9��s��gu���sGr��>�D���k	�����w��f~ox@{z��9�eh��qh;�Q׍�iC#��<����=dC����G��Ф 4Y ̓��Yx�8�y"�}�(E�rM�G�\����=$�o� �N'��͖�ˢ���l��A��d,���d��'c��}��RK��8�-������^���+X�]��I��~�^ό�w�3"�y�����H����F� �ׁ%K��������]HD�ѠG{��~}�e���C�i��~�	�H$v*�i����i�/I�gG�Q�3.�q�~���x¤c�>����m���]d�b�M���~�?����N��U�~��U�~��U�~U����UzW��UfWe�Uɮ*�W�]��W����W%WC��C<-G=��z�������+"�K"�D��D<���/�x\w�0�-�iUd�t�U�pB��,���gyn�7�J���r�\9o3G�tK91�z����8Gd�&����u��]+İ�kVg��[S��Z=U=/�x�燥��c��v]W��/�N��g���^��d����gW���f9w�����~����/������U�����z>]OeU�ͼ*��M�n����l�)�Y�������Z3٦�0�Ŀ�p����g�?9��Z�+c�k�V�O�k9�*��8R�D�h�đ3�#9u[_��D'q��6_��l9��!Er�F�j�X�m'0�<��ټ�-��>�H^�+����OJ$�k�*�[�U����}y��cպ֭6�Un[��\�}����ֱ��F�Vy�/WѾ\�V�j��V�i��}��^v�R�U�\��M�ܶ��}�����]Î_���z��W?�z�)����ktS	+�ʳ�����-���n�{si+��$�܎�N�_kgaG6N���vK�-�L��.�8)��I$��l�m�D6�ʃ�F�<R�[�MR��M"Y�T"[��v�`�-M���j�}��n���2.��sp§CY'�Z;L�D���8�K �gc�Lܪ'�*��:M�M��R4m>'3�smJ'Qg�8NE>������8M���������r_�X���*����/����Z�I�F���V�����_�+��K���q,Dj��/��׿o��BE:mg�H��1%�"1Ok|��852�M1V�R�S��y��X%6�l�d
� E�4�9��IU��^m����v���ɞ��>L������	o��6˼�B�r�6RB]�T+���A����1j����<��]��f�v����F6�B;��4��u:�~@�?��f�E����*����������ާ�v;j�Zu;��}|�����֡$���廼���1WC�X�Giўz5����Gֹ9����j��?d�}C������;{����c��־���wk�<�M�1{��M}���VN�jtرVw�oG�P���Z+�5�7�5+��EL�����V��s���V�L�~܂�醏钛醕��"�+�N?l�[�N�f��[$�LO�������2]]�tM���΄��{�;��t+�-�cn�[V��1ݐv�a+�Rvz�U@�7_�aez��t�������"�[�N?l�$��k�~�8��">�f������"����~�ʇ���*$��w�X�.���p3]�2=���F��e��	�퇻��%o��I��s��y���d���f2(�i��9ъ��\?�iit�;�s9gz�2��M����i����Sz�T�qh0Kfd<�4`Fz~#-U�H���V$��E�k��|����K(R���EQDV`�ZQ���g4di�(--�ِ%��g�4d����*�^+�ӎM0*	��9�9�;��IB��Vf���zi�	fi������8���F:qu�
�����y=��g��Sg������Y�7�ˢ+��he��[Q�a2+͌�!1tN:�����:�O�\h��{�B��֪`4x�a�����d����^��2h�%���i�YRX�R ԵF� �"[�����tA;�ˌr���ò�J�ӊ�(d��\�̤%S��L33��Kq�찬�3�j�4��>�Vg�He�s�G�	�;3�]��1?,+
ۛ�\�"�V�j�
��{��A����\�8:��`x�u��ފ.9�8S������C�y�qY�vJ��V�pP"�oEGjlVXVp(Fpp�{�<����du��me����٭B��������.�y�X�n<^�͏����l��?�>����kCw�G��PK   �V6Z��Y��k |l /   images/7c65d56f-74cd-491d-b8f1-3e526f205bd1.png�W�w\�mlۍ�۶�ƶqc��m6il;il��M����u4����{��RV�B�Ǉ�����������7�lX���������跺³����ȷo�	�&P�l8'i�oߐ��`���߾}�ʈ��{^~xvY�蜢��4,��wR� ���? �TP�����d�0�11o��VY�����Qe&�D�UPQs��fݮ��Ӫ�@	U�����&?���?O�ܟ�m�Z5
�*�C��g�6v�QN���O� }�s�r+����;�� ϻ�>��7*��	�L����<��v��_��`P���w�k[iJ�T���u/�q�(eTulc(d�d�cS(hkZ�T'��o��������l�T���|{Te�/�Jg^��V̯;��-�2N%��m��t_�~�+�N���~|���{~�l�be���B4GZ	���<ߞ�A͠������_�� [����ٻ�U��cL����e-N�{��J����]D�ry[����\�
h��}��Q��#��#�����m��a�g���H`.u�U��/�sG'�Q�������nքY��s�k�mśV'��-�v��.z�?u;_�Q
����͓�r��������s9��Ǜ�s���M�x�ⷯ!��!=����V�׏�o��;��g��-��f�����vxP��t,o��K)��u?O���,�?.��dYqq�$q�*.���9g�_Q��A{N��+f ���Jߍ��g��K�@���'�W�|	J��cM���2���QW�9�+����#�2��ϗk�݆J��.g�?��NY
>�^�x0u0���o��o9h%Sd��-�����x�'X��m`���X��$�������Lz����w&�e�9v��������9w��2��	%K{�!i�c������z�%���������6����hK��V��ACK�(�����p����~���(�������́�hi�(���7�3g#�d�.��
W,t�����q�>��e8���;ބX�Y]]����_��i��D�����������ytĲ"F�}K��myeEf1���g�{&�k�s����>���$V*����T(���;O�|��G.����oV�C��I@�|�-S�����+.t�Ż@��Z]�Lݏ�gO>�Q- �ؤ~c��b��������U(���C��F}��D��}Q���&���E�����1k�7"2an��x�^fݰ,
��1[f��,�=y�m�"����"�ۣ�@M����ӧ�&��܆C�����d.3L��d��+�4��{'�'^w1F��N
�N�Cp�E����뫟��Ȧ������>=0 ��� �b|�2�g��D!#������	yeee��5�u���F���0����2���Y22��[�39#:P��G(�TAk����?\j䀬���P~NO+�N��w��Y�;;�|�I�6�$�Ā!�����kqK��R��r� ���M�ts2��^b=��\U]�o��K�c�E�/Gp�v���N;���'"Ӳ���k�k�nu�r]\\ �����߂�^K����g��5�����__}��f����a۶<6��Q���L,+�����lt��"�޷������N�8b��;C�=�)_i��GGGx��f����a�kQ����5[�^�88�w��";F�R+漰��:2/��OA�mǀ��N��?=�81���<:�Zӷ:='����"#]�=�t�Pu�.�X?F��_0�Q?�Zw����OI�R�z�W<�PѺ@�bsN܇/w�a����y�(�S��q�k:8�0��Ib�������|{#���o�9_���I�2��'�m8�&�F�0uD2l���.\����]j���~�;����f9G����NQ��u�eꎎ^���R�?�ώz�0�S^sYv4�zP�����xs�|���=��.�`{�!��X��dvf�<�j��e+�vN�#�]��if��@����?�,�V�-L�B;5sE��$ZGXq�Ƕ�?��IU�>��;���22e5��N�?uB�\��k�(u�WIC�%�pcYV5�	LO��k;��E�D��p{tl�1��OVX<�_rIog��$�/�d������N�[������ų:�	�H������\�V����Eѱ���l�3�/��U���;�Ξh�z���W�WNzmk��_k����QD�O��'B+��#�e�J+vӤ���2?�mj�=a�~���](�SQ��V�����fe����ZPІ�]9���q��;Ώ7&P�N� �otb����b'4�T���ʀ�.��̕�AM
0d��5,��Q���$i�1�;�)XK�����SR����Ȁ�C� qD���������?Пw�{8)�'��i���Q]���cxƖi���"�6�r����q�Qe�0u-B��NX�V��L�������6e���'��4Q`K���o1�~	X���D��ҖNv�Ha�^�~ex�p<�A|�`���u���3��n�b�����8�O�ҧ"k�7k���`Y���4Y��Pxf6�-%��&G=o��Z���M�'W��%T�6W�
S"�WDsݲ���{���xC��ۭp�Q����W��o�^AW׵�ߊkpB7�n���m�"پ��J@��.���}���Q�nN�<�Sb��b�R1Xk�T���]Y��di��%�j[xVX�Oo�;`�< Hϱ�� �M�>Yߪ�̕�xF �s��"F�k3��&2D��.�ڊe��lWhe�k�$����~�����V����`��w�;�v�Y�E�a�o���X�1]��J%`:�`���6�g���H}���WΥ-��j��!IN��u$I n���?'(-G�@�\@X�L�;r@�� ���2�*��v�w*v��XH���n��ҿ���eg�t���+iŏ�
|)z1��6�? ۔��?��cĚb&�:P�w"r�C�@l�U7ςGE�� ,�����.Z(��gܑ>p���`>�Vt9<eM����s�)>�OQPv������ wc<z��;lζv��q�ܑ.�ܕ�����5hk8����!�'���z�����}d��T
:8�OE����h}�rk�����4d1��k��q'P>0_�pJ�j!�3�����"�����JK���M�����=�P��`����W���fx#4�KP����U(� '��h��I�t=�*l-ksM�n�� �v*���<p����١���s��u�ܛp4�~q�m�e��������p��u��P@��N
cD�gl���/�����僾���Բ��@=v�OUu�jS@b�m���y��#�!>?��!�m��'(�+����l L�h��׆�R�z}D=��2эV����n�-pq���l�K?qP�m����-�;2�qTj��X�ď���{>)<8�u~s��(U�̥�s���#V$)�`7��*��ȍwڒ��I\��v��b}V���H��h$�0�����o��J0�v������y�<J��<��z��
3�T�U>j�E\�QtWA#��u/-N���4�[Y��J�tw��$������H�!�}�(t78{<�r~7
�|���WH/����0�}{�Z0h�����+�Nѓ/�.)��?w�7$K��dDU�:���"CH,��B%�Ր�]J.�<������,�!1�{E�1�;�x��lv��L�8���PC-?nQ�z_�	���?u��g�&�?b�1�Ys�%d�n�Q��1�v)�G��ZΊ-j�`#���f\یjK����3��0�L�ɽ�n��7	�.�R ���}�9|6M΂����@&W�����Q�����3��h���V�5Oy	�+�O\�� �*zٕp�V���y���Vy����>��!��4M�*�}W�"\[m���-���z}���$�����9WO�����]�j��d�g���yU�$~�
>��\�c�� ��t��_����0|n5p]��O¦P_��9�9�
i�$��g�Zzt�.1`70�0R�vZ�!>O����@�S9��:�@|COE`9�m�p���u��_M�O���	���)�����q<�y���ᐊ���2���QY���u��0�.��"�i?����[Z�]09|���+D�TC�J�B9,+<�c�|�e��
҇��V������Zh�s/����79�b�_I���@�k;�*��q��]��v��n���_)����Zi	%3��GTSF9H������K����ҵ���4��ޕ�AQ�7���T�;����z�P:!|frs~J̾ W�-��w��4�{q��~ �����J�C����[��� 2�fk����
N|/�h>����o�W�6t"�)=:�o��r�p�����Ts�핂`��K�h������I���[��/uY�I�֖1� �9R��xJ����P�;\ju����yǉ�,|��UA�-֑��q�RؘeV��9w[��NW�Qq)��mj?�(�ʏ��cBb/r)�jl�笄�
NSPv1�[�a�P��7{�ùam�(k*��h�q^#��T���ף#�f�GN*Lk�]ǯ�-�q�H˞SfÝ��m \+G?�9�v���Ep49#9XT@z��'5ٗ�
�[H�*��>nQ��ܛ��em�&���tJt����f��b��FT��<���b82!4M�yD��H`Y�A�#�f�K:����0/^Y!,��0�]J����,���e#��N�Cy�(<�I]�`���$㳅(����]�N�����m�?�R�=}Q=�U�
.����;���HF�\^s��Qa�����u�������,�M�MC�ȗH�^+bP��a�E���Y���=D���M�M�e���݇c�??�WV�_dፊ�C�$�N��^�jۮ�t�5$T�f�6T�\�5~�G����'�Ջ8��d���~�d�v��5D��^1, ��@S��V�N&^�~F*�bM����)j�.�DE�xVy���T9-c�q��s�WGi?\��}5F�5v�Mf�eV"w�ח�?��Ki>���\)τ?$��#�k�x�&���F�_+��}��b2�D�7����X��1O��0�<�-���$�Ǫ[^�l��A\�m�]���.utLg'�sk��:�ըmű+���(bz3:B�ۈq�82wm��<p2�$�ӉDvmr�)ɋ�pPv`iu�MXc�I]7e�ч�=��8�h�=�7�N�`ɠ$E�� ���{��E�{0�mPO�`o�t�4��c����C�b�܍CL6ɞ��0rWq|zQ����b�e�[n�h`�'wU)�����t�fX.؃}Zt���ⴷ*�D+Q��NT*�F�'Zܚ��Co�	��Q���`MZ_�>���|��2�����Q�H<�[���C�@����,�*4��_k�<'����Q�6g`�wx�*ɰm����@�MӴi+��K�J��Y��G�%Q�,뉚[��F��Q@Gǩ�h\+V���]�����r"`e����|#y��}�$��8��E����qJ&>��
͑�.T^�(n*��>����>��G�!A�c��R�s�O��9o�z�PIe�qn���y�K������^�Pa�����}�i]Y6�)$��1�I^)8��~�p`i��++"@o{�"���@g��$�����u�h��Z��M�[� g|N�?����bVg�m]�tٕ���r�:G�巇�:Na��e�!��6}�D=MHZe�[5��Puqa�{,���F)u� �4�SkT&�7K�����rbud�Щ3�kpbqb�C�E��L�;���Հ�n�	CĆ
)�l���
�[s�Ϟ�p%8�
3��N&䐃m3:�ћp��*����h�h���ڕtXjt��UT���+��}��Rg��dy���`�ڡ�\�&���j�TKO�7TVGc�,��9R\��2lbGPi����!mʪv@m���BE�����ņ�Y�0`GY>��bΙ�l���+�w�B�h
E�����;�LU�%z�[ں�1�܁pP�s�1P8�G�g.�a,.�'�ZSQqٟ�mU;�()V�S	3;U-�8-/�8'�6n\)g"�Z!�U��9h�*�h�%(n;=2�Ť.!��	kZI)j�i��	�M3�L��J��?V���!�P{��
4�3�b�T���eq��8���:��	j��rH��Jه�Ĕ��L����l���=u�) �c�*��0��T�:[�Ɋ����Q$Q���Q�$�X	�N(I������Wޫ����N(�V�*�L����%o���觑��.�� �q�i�zBCu`�{��b������.���L�؝�<�BmZ~W�?�G8}'��7H�������^s)%�,�_��@b�}7Y�S��;� �ڸ+@NE�m����[�Էr"E��p]_�Mϰ3_�l'+g+B�y�X�z��Z�.�V���=��<Š����*J��B'��v�����]1ԸFu;�%\?��%` o��]=h�
j�yu��:r��]G���kqN�<��R^NJ#�Oz�՜$�2����FC���@���+�s��AK�
t� ���\_��6ݫ�.*T�e��~ps�lz��(�Η�O�L5�A�.�
ň$On3Z���Ō�y��u��^aXqdS����&�������+>XY(�w�Ale~�{�p a���l�ks
�UĶ:��u�Զ�����v���2"��F�q�YSڱ^%tc�b\�c��+���}}N���xɘ�4,<,���Vh���0mߜ�b�}u�6�+ky1�왤���~����_�b�#���\��ay�E��Y����������4rR�m�C~�˨�1^��]ш��d���D�7q����9]��~n	��%T��`���))Ҫ��C+�s㈙!���2S�auԋ%��JN��0���X3��������m,�ٲxYN��@�ՊKѿn6�"����j� YF18M\~���'a)�Ub�g�+X٭��Q��z�ߌ�K��ͷcf�_�X���\]���u��H����G�i�H�^�����2�;�L̅ŏ�?E��C��һ��̶����ж��i��u[��>��Sp��K

��+�(��W�T�N;�w-=|d���!�&���]Ʃ�������-\�$5��6(?�[����p��AҎ�?e�4�H��sO�LcVs�H5:H��Bd6[ӆ-�.0�q�a�ص��ﹱG��+bDvu�9+��~g�qRh�RBB��ͩ��ҷt��P�QW��Κ>�j��MG�S�5�GvΖʬ#*���u����x��������檥B���4.EIW��h_�&�B�w|�Q�l�z��U��Gr눍�hJl^��]k���!�S�*"�]�8�i��}�.�Fiq�,X?/-�/�=(]��,qu�	?��B#���_��Of"҂�]Zj�Ԋ��Ɩ�U�!Afl���'%��Ɖ|�>�c"%߼^`�HZ[qԜ���Ȼ(	a$�=��U��W�������lk��P[�Y��{^���(���>T*3+:�*,���OֳG��[������b@��t�!�o�E��'�"�'M��.����Q��%��HkUk�
o���A��]㩷C���}mIk��$��e�$�<�XF���*�5��DxL��?AF`�3�*h?��PI�,�P��.cR���Gm��.`��AؽeEl�bFSw���RGg>��a���"ɣO/T�{Ef��>��d��:�*����
�U��:������Qj MW3큛���8-��>%)���-��t�M���H�����;15O,��^�_�=���������.:U�n`�
ܧ T$Z�&��4�r�㥨ܺ�>.�O���[���9ssi�d.n�7�X���ȑ)��dXh)�A��J�U�Yk����O�+(\h9o��������-e
�^W؛�?��WE~�����}������_��
=3��t|4R�Rm�g`J��'��c0� t��zoS��dz��R���?�4D��M(d?Ǆ�"��0S�8t�z�.v>>���0�X'|������y�{
%S���D[�8�*��=�f��[��%FJc���07���IgYi ��G(�^BY����On���)�b����ͼ��rn��;&_�$C��.�pi��a����*�K~]D���4�Z���d����Y�/�xȎ-��*Bx+z����Y
e�Qie,Y\:D�2��IBF
�Đ�@�<k:4���������`� D/l���񡥎����f�k0��06x�XC��"��m�6��>��Z(^4ny����	�H&T�}����j�pI�d��j-%���iDY�U���7ޘB���{�N���M(����=	Ǎ|9:�C��Y���zDJ$+�ա�¥cEj1�d�&�[�l��HL;�T���I:-��� /�C�m\0pKa�:��Mt������к�?��zD��Q�L��G������o�J ��=%N�A�w�WE������ơ��x�t��jeB�EVs����P�x�-2�kP���B��ԛ�G�]�,�f���5W<�n��(��+d-X���h��vpǦ�͡�eH��j)Pv�VP��N�~�위�aF��\��ʖ������{���6��AK@�؆a]��(;a*o`��U~{�|���7�h��5)�)roAeN��W+����5�ZN��%>sGr0�T6���=R�l�.�7����R�*N	ș5b=�1�=n�2<���ᷕ�t�$gl���������sG.��s�����S��<�w� )�����w�����1�U�#@w����a[l�*�**��V9֭ߔM�5�[�q�*��4���]�����	��]��$Gm�'�]녦�Ma�^2��^.�:ص���
�V�fFpF1���ٓD�+��m�_�,=��ZP�Ga9[���%�L �_K�Ѩ�q�3�<�%��{���%��ʩ�w���p)�qbJ�D�=� H���mn�}���������i8H��/�?t����ˬJѕ��B�¤ŲN���`Lh9H�q��5���a����m� ���ޗV�ɕ�D���e���	�� �u��
�h,SZ�%^TT�S�n��Nhzҍ��B��y������~pH��ɉw{���C5Ki������hύ���@��� Z(Ejsh2�AL�~�~���I��m�U�:�T���5fA@��'��y�~����1�k'\��k����0�=Ǥ�97�T���b+Vb+���W�Y�Qr]�r��r�:�DF�[�rr��*�W���ET"����8-���|���k���*p7��y�>�lnvo��ڵo�l�u�=WQ����.qpGeG��t9wJ���x�m�P����Ӵ�[m@��Y J=36�-�]�M�y���o�P�"��s��'~�n�u�Y"Z���R���/���[�CsR1�*-Z��
ݷ�xqr_���$i}�ʙa[D1���r���+G��'�;��
���<�.;�R���kCy}<@L�/�dk�O��6�B��{	�3��u�S�CO�5T��+�683Y$�!r�[C�/!�jG)Ţ۪y����Q*�F��ui�����K
|���$ph�����5�}fR�6��Z��#R�h�0��wM���9pm'�2����h{���Y,C
#?6z#$hϓ<%����tn��,x�l���Ѐ�s�)7Ke[r��;i3z��~G�7�a&�x���'����A@`�1$�;���KZnơ��I����k���W`� GgKXz�!�e����h��ܨj#�W��&"ت��H�p�*�>ƫ��!�<�5d��>��n���5�����Q��z	)\����`�=�9꞉`]aG�O�]��<	<(��:���K��I���)渇�!"�?N�a�_ѷ�]�M�f��>ux�2t#Ƞ����h&��?��{�A"*��cs�'�"���1m}̷�Z�����?V��;����A� ���w����1��x��m�h�Nq�ki�-�Wa�ȑ���2�eҲ���0+X� ��-���7��)����W���Ɍ�l��fK��A����f�ಚ2����B�z���JeW'zF���d��p�d�){��n#���"�2�	��g�Ӵ�0���h���+��C��?7��9��M��XW�����t�����|�������'Nj���Ӱq�F������Q��#w���靿\��gHC��_�r����9 ��N������w�
(vN�v�"\[u��L��5��=�ט�5R9��T�����i�3��k��`=>0�%_�	����Ս�!�ۉE\)3�ֵ伇���I���:����\�i���{�?Z~ψ
�M�靖r��_ʡ"�B�&���k�
6�.�f8����,i�I�v��Q(!I$��%�ȩ!2�Dځ�B�{�\���tohD���9eM��y�ƦL�?��7f���3�'�{-��1���U���+�,u�@�^�#zaּ�`�#�ňћ` C$`����3v��d�t��l���%!�;����I�:�ћl4I�B������d�[��7Q��ɝ�jj8;�f�)�z�F�w��1�$o�{�lW��Np4�b��Ζ�|z�WS��E4�J�&^n�_��n/Z۫�G_��:�f� ���C�Y�GЙ��f�2���Ӭf;���]�$�����-��|vxˆM�F��ӊ?# >�#��9��j����4ws�z�$���G%�
W�#�U�?��� t�����]�9�֬^�����<e~���ˍa�ʶ��I�k��eэ��Ki|��N��\��MC��BԐD��D���ToN���U4����me�@E�Z6u��$���%3<�ok��R��w�������~b��?-�Ʀ��Q�^B�3���xh-�z��>���)Á�Wt��ŝ�ُӔ�`��÷2O�*�lT`'h'�YY�iV����4�I��Ĉ,YM�Nh8�	����7oNgXs^۟\5uI��m�U�;�e�K�	4~$�F��H���8�~�"�����Gz��GR'�K[���������pA�x\������M����T�7� R�F�0;�So�%ݿ�G�N�%o#~��_":��`��,?ɪ�6�bj�p`>��X_+�������l�B	�E��]��0��I�4��*2���a������F���Pն7�W�"�O��9`�sQ#j�XK�{<��^B����M9v��{���q~b���n|]oq7G�CT�#�Ow���vgƅ�wf���5��>Q����hu�`X��_�&�vW�8�r�W�����jG�����y5����p��ݮ0V�&��s�^	�\����VYN����>^c�����r&V[_�p(s��{�
00�.2�+V���	k������j���A��ŋ�Bs~����u�HO;"F0cRl�����i0-v�r���"�+ x=P*?�W�7��W?X�?C>�U�5:L�C0�ْ\�ˀ��ٓ�ۛ\�vʢ�/.b�b��t�l�#p�|.ؒ�C�k�{��������� u؆F�+J�F��������W8"P�"�B�$���؇H1J�~"�0�.��r}h�X�7b)����pSТ�_?�]�V*� �B�c�{T����ȃ}zKtX�t���V�a	D"?�`� f��n��+߬�S��|rc�j�U����D����.E�>�Zz���~��@���-,nTճ��y�p���zMks��
�AVU��*pa7KY�l�蔢�-0gt{A�ۙ�(?#������n>^��e��R�ǯ*3�� ��`;�q��Q_A��E¯Vc�ˢ��ǅ="��~�c`W�ؕ��)��)�+;M�	��^�)_��i~�͟A;)(�� �}R����d9P���@�B�ł,�*���;�]p��"��{� ��.��z�i\\�c���,\|��9���2|R�tC���8ښ���-9�D�ˀ>���^of�����/iB��	�"8-��.�����=�͏�L�����g$
@�-���iJ!��m{��4��m����F��7��
���Rxf�@��&�YC�i'��}џzuoK�9�k�8�p]�k �`�@ɗf���7�ݽ%�Hr�!��޴��a�k�HI�C�~�C�ְ}8�	8	��;w��"�z+��c_�	AM& �+ɂ���@��C=�&��h
I�[�-�DYY���hբoW��h���<J=��i'o�A����?��Q� ̏c�/��w�Zǯ��v�x�O�dC����w?���m �o�Kv�����b(��+��a�/湧V�a ,�1jY)e��F*���쯐�V�t�������V�'�`Q_��i�\3����T(R
֚\������Y�C����C��Cl�a4��N���*�3�������1��JI՝���V�8���U>;BT'�nj�*^���d1[����d�%�0^s��8�i�FlD$��y3N��?tK&k˯�vѓ��Zű��b#�P��� Q¡$�߂V���� Zϙ�|`-��B0��.�hw�2�=a�����T���w~�p���8x�=>"���}ΡZn�_�uP���+�G��ŵo�B.U��G�U���y�Z��O��"M����'	�!	�R;�1�σ2�d}��� �7b�k����9�R:�N������A�<(� �S���|rn!��^��'��	S�)����N;��2�<�G3�x����kWta�E���,�-͞ �/�ұ�kr׌���-�.{vE�%ۯ��%��Et���e�i�N�)��nD�j�9�n�5ت�A7����'��4���8��0�k_�p��8�q+����X����:Bن�NǀCZ-�=z�d�����r�Jd�0O�)p$����.�FQ����MM���dۀ�����	�0W!����Y����'1�-��(3�2�.*���W7}F���~�ż��@��<^�.�a�O��Z�$'0Ӥ�Pw�}ڻ����R�Q��r����e�"�(�z�+�S*��Vۓ�����+��?��tS��FM-�!o:�p���u~�>+^I*EJxi�v�Bb���J��ந�Pjm�iCi��^
Z-��R�����5�NI�H�}z���	��c��Uh	i�ʠ���t��ak�hg?�Ӑ�(���ҊSJH߄�.��|��%��?k��҅56��ۍ "u�Y��s7N���bɐ���>	��J���?�ut���{^
o||��^���y�;~]]^���{H�
NY����!D!��˓]|ۖC
��N)Tv�7�z�$�z�����*����Q۱Gn#7��I����0���;K�1Ev���FG���"O�n�m�8����T���>q���R3� Y�Y��Ao2�aw�����o��$1^����}�0��2��ּdU큗�פ8k�͍�?$�t�����5�bv��['�Ɣ�_��n��������`n1�,|u`����( `y�CD�Pm�����
�o��W��]�?�O+.,� ?�II�v�5z�f�.b8]w��(��ؓx����#�D����]1A��d_��|�k�'�'ۄfa��.;%S������Έ�P�^� )��OA���"YAE�!3>�˿�j���2""e�Ҽڛ$��P2zu�p��u�&d1����o
�L�J��B���8��,P		7d-�v���2]Q�]o�s�{�a=!��w��HO�P'����>��"�&����C��Y�E�ť|���A^�9���l_���ժ��
f]�9B�K�|�I�19x%�*�!�.8���ѡ���!�[��T����4XT�����z��M�YH+��LmoPAt���#d��R�n``�a�B+4�B�t�o�yU�*'X��W{�R�^4қۛ�G����=��~�����o}�hucWV�-�=Kdi����o���9٦t�}��em��G���Q�Cuo/)�"I���	G���߶�î9�	�~;�<�}���d���O8��9����Fg�z�w=�1.G1։�];�ӎό�ŏ�$@Aſ!l��0�MS�� @����o��[�B��Up�LO�Ž�4�2߼���xg!S�L��	�+^�����8���.�v�m�SPC��Ё}� f���E��C��fқz8��CV}V�W�� ����H�h��R���`���)8���ƙ�p���k,���嶺(����؍,�(3��G'!��	���	������v�X���9���ڎhź�k6��8�l2世V꒥Ei�\2! ��d�X_]�Vm��D�"�"�?V�,��s��S?V�p��e���n۾�?p�@>/Ch^;ӷ��{�{ej��٢�󩈋2g �JF���,I~�=o���DKm��2��2��hU���N��v��~Q�j�P#<�*%%�ɉ�Y�ߴ�[	�t~l2ܱ���~^2��Ň�8��w 4h�o!~x
��2`���=�
5�lڳ��n��!��J�/T/`Uo��ư�"����/����9�*O�N��KU��W��@\zH�g
�i_:�>:��L����UXa����y{#���iX�S��;_
/BG`����n*T"��Z����I*b�怸��V��]�
�
]�p�*��j�t"=�~��=dB�Oܖ����7}/�K�V�5s�3�,��)��٣f���c�Vo�~���Aj�P6+��r��*C�w��983�ԪI��?�"�)V�u���w�%y�G$a�P.�j�z�p��a<�nۢ܅F������'4�f�R�{�+���S��'��||�p���DH��P6�5+�WQ��u�y˚w����.&�I��*ޖ�Paߨak=�����#~N�aJ����d�6����n��+���d��a�6A-}Џ��u�rZ.8t�u��8i2r�}��&���s-�+��?א�x�W��,��PD-9�g��&w ���#�t���yW#^k�������V=�ά��J�g���M�˭?�-��Q��i�rV�e�m�g�q���u��O����^�����PN��HZM�6�r���^�c!g,p
x���(ml1��V��S�3*]@>�g�"�1����)�e�
�jp\�]�f_R�3#��o����)���Q���\rm����V�W��ȿ�4a��ɪW��z(�i��HY��h%)q-D��1/ ���a�p������n�Y(�
˜�Ʈ�@J�y��]i�*�H8(�T�j��їĒ��	��eA
���M��V<��5�$HZ��j���z�{s��:�S�:z�{`�#�߫���QN7�%�%N0OЪ��M�.�m�o�)��V�X�2�.�����-�:�K����:̓�����l1�M�\߲�V�o`:)EuC�(fɣO7���m&**|ؐ��)f��lᖁ�#rbP@�C�}'r)A�3��qI|�pHx�V�{R����U���XC�f�'S����Bs�|&Z��W*֛��|�3��"�p.��%7�	+W�+B�\�R&��bEѻse(�*/�jʗ�px*���|�K/��VHƶ�A�Y�m�����ȧ��h�ô_��6�zx��X��P"��sp��MM�BtӨP2��?�xk�L9��Es��"j�
@C����R����V㮉w�D�2�)hD��"R�;�>	���lXc+���@���I<���Ռ����,�u��nؖ�b�.jM7��埿����(%���v�9l ��&	xeX�#�,e��Ud���f(���i��4�1f��7Z��J0^*�y^���_�!�إ�����n5�h4
g˷�68�`w���V�cz
��uH�V;���4�ߪ'�G���	�Sm�a�T{Y�����l*w_
Mvb� O7;Y�_h��p$Jc��_�E�"���ی�I�QC�-x�[t��"C���#�&~����?.
�\��&��2��(�*��C_�JaӒ�S��Z�pc��Ҩ���M�n��#�M���`h���Dr��~K��R]46�F}ޓ��fpbo�4���5I��xm�n�<�n��!Z@��P�4���ʦf�TA�� q�p�0 #kI#(^�����%��r�	Dq[B���~󦇩�UqhWPo0��2�6���������WH��-B*��l�\�]� �.���/�J�0�``?���e�F��,��:�)������Ԋ�	3mY�ĳ��
E�}��|�5@ʿlQ#4UIUL��z�yJ-�V�טd�ɮ��[T(����|��$P�:0H����[�����e �u8WǪuN">6�m�\�
�Vpx��Q��E�F����)�5��%><l�v<�,Ȗ�fOH{�*0�v����C�k����I[�48��|�l <�ŴnN`s�	��0��I��4Pa��R�,'��W3m"�=��-�༢����#����jC[Rt|>���1���`a!#K3\��&L�t���"������lNk�=:�e�KK��	�a��e�q�F�ȼ��LX�0�Z����}�h�P[�[����;G�Y;9�����N�^bWά�A��:�X���0*�i�%����P��bF���|h�$�T�M*���,�ܷ�ؑ@���]�s�x§[
1��=!�k}���
�j��Cl������i�$���{�;|��]C�u������Q��6�mB���;��x��q��x=ś*��Ɓ�m�8��脤`e�1IXą,�;�d��1�UEU;�^����2��U���#M�C��h���,ʥ(�".ŉ�y��*$����x���/��>2 :6ER�U��"s�����l��b-I�Kb3�F#�鵒�`����Ӗ�I������QU�$�@z�2K 2�
��Ј�N��ĳ��H���.����i��:l:E5A�E�7�Z~�@ӄ��躆�F���c$���D����r���Ǵ��!Kl�aCh�%:(�a�\�!�9�1V�������{�Ȏ�#�B�.��98Kr��MK�e���5^B��HR"�r���P#��K���z:��ȴPO�T�1�פ��i,���G���PDY�(5F�qP!!�ns>	s��Ю�6֕�`��+��0�b��&RM�X�R�L�LG#�x��tHMC�+�*It����B+F�@J�T(iо
��}P��h~KK��	�OQ�!��0�X���֪�Pn�������ǽ��!}ND"C-Q����i{��$V�%�� R��B��G�±�Yh!��h	(>��I�w� ��kRᴥ2kc���DSj*�'�I���~�~��S�q#8k����%Y�ѩp4���	0��I��<a�<�D3J5��2N4�D1I4S��1��5�]+rf��=������ĩCo:�VUw�$Q��5]��nJ������7����q�j�x��p��p��h�v�'�'�L�kL�u�rHU)�u&�U&�3�:�t������b��X��X��eӜ��ܭ8u�'8v��ߝc�b�	�s%&3POQ*d�H�IZt������S�b3�$-�tݔ�/H�!j����ө't�	2Ze�v79�/n��(�Ǡ<�����A��М���YC5k�l@���7��$��Cq��:�b�b�~��\a��@<I�6PR�ٳ@j�k���3�lC?_MX=s����P(8Z��Wa��tCW;:�ѱઊzR�P��qC|�Nf&h6�j��@�!3<j��lRnax�F�F�L��U�a��$Q���b��Ү]8� �Y/=���)�"Pu�]�i���D�/��Kl��o���p�%ʴO�������ǉ�0VU��u��HYo4c�1ɻ4��r4��}��^�F�ˑ�⨯)��)���{OQ`�!I4Y�Q�K%_v�:u���`zFq�e�q�u�Eǫ_�\{�@`q� ڰ�9�3��b��E����D�}�8w�����v�0S�����풊�uv:BTb��J��3g����b�SGo����_�P~�JXI2^�$���y�y�[��?}�����N��&9I�	�#	��"s6#ׄ��V�����mh2U���B��*2�x?f�RBV��f�Dל9q���S\���S��K���������_���X\��9����#�N������l4Kh��u�I��<	6əL�������i����Ҽ�%Xb����*6��4Sa׮=d�.���~�v��Q��K.�Y��(�<{{P���i�%�x�7=�yݟ��w�����G����c˚�˻��r6�V7װi�����к+���H�>k]��p�~��1X����6��dХ;�㪆��L�p�������_�i^�K?�K�ehi��0$X����t��d�i��`G=y�����ݾ�6����]���=�~ͫx�3��Ն�hXX\dcs�?�����Bc�O_�~5_��l���	շ���Y��u�>
����ٳ��hL1q���|�c�qr�������׽�n6pe��1Y���<囿����6Nn6��mP�$$I�R��{�4,���-��S����򎰵Ͽ��+���p�AגEצ<���p�E����c�`��*�݌���r����-�����ﺎ�}�z>���3�6,�>@i7u�NJ�A��@�37��T��gӲ��]-���*q
mS��@Uy�a4.8s�$�W���=|�c��>�B^�����[&�E.���+.��bN�ӻ���{n��&Y�]���&aZO�&�)�X�W;{��b��ٌ{F�s�C����y%TR�RԵ��ѵp�%���}K�z8�|˛�՗�����,�HŴ*�������@O�>�����bQ&X^%��7|��5�����gPׂ����z}ֆc���o}3Ֆp��h���z7A�d����nrk��W����ϧ�@5�C���2�L�X޷����_��g<�)�����[T4^&D4�~o�1�U�mPZz���r��"Ck��
|�{��� /|��r�'?����B�8L�e8-X޳�_�����o�g⽈F��*(�pO�nJǭ��-���?����v�f:�^/|���Ka�����^v�j:"��X�2ٜ�%	u1e��2������@o.\7P�AB��v��r������Oj��\�ǣt��L&�V�|ړ���[Ѣt4�)"B�<����z����+g�ҡ&�_~	�_�Y��׼��<�Ϥ���W�G!͈u�]\�[�vmha�Ǻ�IO�K"F� \����׍���<I9q����8r�z��F���>z}��:������K�(���w�����E�A�QTu1{ڢ��]�Vo���/�����sۢXQ��ህ�%��t�]N;ɧ>����N;� _���(�$�aR9�ɩ]����"�������\�C�0R\A�C[C��p8��A�EE?����Zu\��H���NB����I��nP�,���?u�y��x�k��S�O��!�-�X��`e'Ϝ �	_���>��˻��ǌ6�ƪP�^����
�0m�ͤ�Z�퍸#�c�1P��(/�۽�=K+�>�ƿ��}��#f���h�SX�J�{9��!
��w/���Ե�J)|0rQ$P��/_�j����d��0�L�{=��)�{VX�8�4�-���>���wf]���ըv'8�w�@GbPY��RB��
�صk�z:A�ǒ2-J�VV8�z��^�mG�K�J�&�����5:���8�So�����Ý�����0`��"��L�c�+طw/�����_d8:C��2�4��t�F�!HӔɤ`:)CH�
�׳�a�e�%H�Ci�wu�&�1ܐ[q6(֣���6dV��UY������P5�~g��pD�4(l�a���k�� �IIm¸��"�8��%�<�S�'�������ޒ,��������X(Ej\]�*Mb-�"����;�Ž��㘷����g��@���3�LILF�v8p�!�N�F{8xhO|us�"�vw�-g�Ӹ3Tޡ�C{G5#uA��Q)l�6(Ǥt�$Ǒ �����jE���t�h�.�)�NL_kPVϡh,ʚ�ps�9D73Tq���t@�P���(4Z��ZW��0�N!Q�!���F1�Kl�Kwi��՜Y[e:a����,XySUbu��5Z�쌙�p�����sOe�5�
Lqv��S�
����[��Ʉ�搪�I0I�N4I�JS�#�v��0@UNO�Ԯ"���!�q9a�F�L	��T7T���CQ��Mst�"&�%��	&��":�EE�tC�CϘ{
;=�lN&��L
�x< ٽ{7�k��C�$#1��GN�/Gs���l'<۱b'��m���wD-�DB�H��%��r�AQQ�N��N`s<bie�gN��-0��Z(��+�$�$�8���&�|�����,��%��F=�a�7�jC/]�&���@��7YZY�p�d
�l��u�d8��LA���Џ���R#�D�D|	>�[�M�#��E��v���2b�;p�w!�)S	V)��d6vaw5L&%h�x:��2��fZN�hև@Py�q;EY0.&�xt�Rᨼ�q�������,�ܭTlRu'�����S�J,��)�ҕQ����C�%�eŤ
L�7�߹����""�{��09��X�\������8��Wu���N��o��|ĥ`Tt��%AB!+�4FL�ގA��³��c]dZ3�)�1���R�<��������Q�����IM���ׄ�)��5$�FN=�[A�(	�FuD�`g�bM�V6T�ߎF�����R�iC���yJU�M�M��&(�dZ b�&Ӑ���$t�ւՂ�=.�
A�U����[Z���|H��H��LƐ�����V�w*�5U9$O4�L�Z�*�U��V�ut�и��,CDpN�2�4:�����l��6�:t�6oB}'����υ�kJiA,8ݐ�	�j2kH����$��]5��i����&t�ݑ�>/�KWP��Y����^'��^�O�w��)����+j�1��Ř�&���<vB�C�i@��w@/>"sGĳ<�͘�`i�^����<�=t1�A�4uEb��(��4M��!#M:yN�X��)�I�5��YG��j|��k?�&�k��E2���q2����xUYP�n���2M�ʒ�+�ص�_y�2H2�+��&KS�ֈ�4�	!�JaL���]�2�m$�Ѥ�`��h�6�;G��6��考�&�%�"KR�������Y��(�(�#|U��;$I¤��<�����WUS���.�s���G\��v�0|�ڿυ[1��{�*�t<E5�L[TR������I��P�z[:�=��2�����9d{k�&SGjsƓ)>6'k�`i�"Z�D@p�_+Wۜ�y� E�6��[�LJ��6���pL��(��Ťb�����c�C�\��좚N�W,-t�4R�h|I�L�C�jD��~�8�mGL�[n���0j#އ8����r6�4���T�����g10<����&��tlJ'K�ur��]���F��,뒤]���Q�๨�xl_�cӀk�q���c���ؾ�u�}��d�zz�����S��t�����:�Fь��mB.���i5	]ڵ���xW��r�e�M�݌Z��ݭ�d	�����
R;#��2:��q����ۅ�`k;�21$*G��Tn~'s�`GUJɎū��6�B�h���(�)�^zӲF��ӫx����!,��ѷp��K�"
���N�sB��p7?h�fG#$����<m���X����P������3A+��&���Ӑ������6��]��	&v�g9#LҲ�~���N��@���Q��U����J�YlhC�ky�r�4\��M�)��$	��~�(ʺ���JG#��Qk�
���h{�����䨻�J`s\2,��4��EC���.B�_5�$�(˚ť]T�a:i֡���jZ`����!���g�D��	�w\�g�v�J{��$I�����*e��S75�@�!�R<�i|0��p.7��8���F���貫���O�(��W�����oGK�W��2n��ӡ����ʀ�?�qۮ<�$��f	2�lh%l8O�1:k����|Uy�v-s���˹��Y?u�z���X[�*����(ȣ��
�w�lN���<�a������b�"O]�6	����8�CL��	��Ϙ9�6�1�{8������{8q�8���q���Q�Bj-�I�y�aay��x��p�G��'���S64�7����p��\DGQ���Ϸ��%:Z�tcuo�Pd���0��Y,�9�ī*�YΒ�:ư������x(_|�Uh�0�B�Ȳ�N�C��`ƊkH���ĥ���	�l��;�(Oє$V���j�o<&��~�o{�?��5`���tJ�A�t�.g&k�������rN������'�K.���^�E��~׵�T�a2���C��,.s��U���^�X�3؉d���mf���R]gNm��7������k	i`{�Y=�ƁK��/��|�s���h5i⸽���������|<FS�,�Y�ȁ�}����/x���W�W�6��J��>t!o�۷��{{��&3�ze�aC�;B��S;�׻��6K�j�J�U��/��?K1�Di����M@2R�R�S.ؽ��}��XY�NC��F ��P�,0�v!Iv���Xw
皟�uV���8�+���.��7��O�.n:|U�!�	xO����7A}�4;�N\x�Qc��ҫ���Oa����g}�w3)C�V�h��S8��Q^�ڛ�X�{���8ҺκI�,E��gKX}�1��Ϳ�J��f�=L'5��'��E��UK�F����|��u��[�vq��ٟ��O�:��ޒ��0M(�/j[S�mOw�$1�cu;��`�vB=����A/a��1_���=�/�N[��W^�+�h���PI������A���	W=�*
�rUAYm�����C�L>���r�v;�{���B�@?I0���əLk�����Ʌ����J��� '��w������GYLrV�Re(����CI�8F5_bTB�PT����N� ƴ�GQT����5��c��p�/$��>�?��?�7_��|��7���Ŕ,OO'h�=T8'�^p����:�C��\�g���\��g *&-O6ٵ����6����O8Q^B�v���Q's�`���a���畧tM�&��J&��U^���sG�g!�z�$y�eq`9s�����~�Ϯ.�:�r�SD,�x�������u~���bbv��~�`t&���mS5v��,�t�e��v{l��cd�b�`��j�'<�2��)��'^�����@�9ay�^�Μf���<�_��������=�ϔ�<y�`qq���J���m�9b�m���#�#�,�B]MX=z��vx�W?�o������_��G��6f��]������į㍯y����ȿ��n:̲IY�)��1J�$�}}���`��Z�.�����ܑW:�	���4�57m�ѹ�B��ky�K^ĳ��L^����+�yƴ(!��e��|abqO�8q́���km�����.斛oW�}-������"��8����>x��}�r��P��g�ܤ��6�3�7{���j��Z�%I049G�4X
R��� 1i��W��K6H�v��a�y�w|)_�/���/��V�׿��<�q��ſ�&>�zSs֦hk�����X�$�~�Q��QT^B%@u���1@a{�����E�k�LI)�׏�W�XJ���t��W��K/ Qu�{\~%�����3%?���D����A���@DBɐv?�y5��#Q�ukA�ZBs�W�
O�k4�/�M刬���]�oy�y£qš��:v*��$�C�}/W�ǯ=����5�N��5�,���R<N��T�h���ǝ}�ς��w �b�P+a�a=Q�I�t2~����'o��?⫨Q�¤	���:'��y^N��|�O�v��:x�ë�֫p�!F�(beu��unÀ�E���t�W���é�r���GlLw�h��b��;x�ATN-i(�h�����>��C��mG�t���:I�m�F�ԦK�:8��>aA��e��HX������.Nu�tit7�I�p����:�U�t��� � 1�`�׽���wv���>�,�l�ڦT&�2]*ӥ�=�ëQA�R	FE�SܿN'�e��J�Ʃ��z��G5�{�ڷ�z��;C��Q�=Tz7��M�v�����^*��X�}j��GiP'�h�Cf�j��iJ��	� v(��(U�L蹆ASӫ+�����ꀃ�aP�Ϫ�^�n���&�@��b��ω��f�T,T%U�bS��T,�����~w$��P+�ހ	T�="Ģ�k�"!���#�C�<B����:v�
h���B�c=��X_գ��&�,�$)w��)dST:A%��p.�����C�H%�ڃ�Q�No�mc�O�tR�b��W�KE�1d-Yj�&��:Vȍ'�B��\k:Z�1��6�C�*r*�����	�K�Q(c��|�������ڢT��R��btM'b��9�tѶ������ִ�aM��p��s��=�h� �W��>|z�Z�eT-�>��^BΩ=s��*��C�X5Hw�P���6<7ي[k�8�h:�sb��N�煾x���6��g�ݶ�T�s�~/������,=w��?�
j5aA':��
۪P��Ɛ�6k�Q)�K�R���Њ>�V���|��c�S�:�3�M�ߖ�EI�N��P&J�`�ic2���g�C�WP�g�̇'��V������D��5
k��u{����Z����ʦt�C�U��oBd�V�D�@�އsM����l�D��6m�/[�dv�6!��S:�Va_���vBe�w��4J��`}�]��G�dA�����t�ה���U�v
b�c�#~�d�5cH�������FlC���XO"T��2�CJK#��_ �袺C���;(W�CX�am�l��zD�C3�mp��u�X�XKc4�cq6�5РE-�
�a-
ׄ��VG�+|#!w{�qj�8��Z��}�C%t%a���Qa"S�(�bV2��
6����Ah�Z��!5>&{�����b����.� �.D��c݀!C�q9�w���Bw�%S4"a��|\���
M��
���ǢYM,�0�l�^��Q8+��m�r8#�1�=7΂7B��@�
Ĥ�$C���qw6#�;$xRj����mMܺ���e��`s/�cP|��Aۓm���e=Dv�%Q+�d^��,uRI�
�;ʮ��"�-h�6D#�oڄ�s���	!�
��g瘠ۛnHH�h�I�ǭ��7Eb����)˒�	U�mbx��$4du�ȳ��R!`��3>TT�!Z�#�j��-j���c�!��Ј�I�N�8i(����R7%u]Ͱq����D�����.��B%s�bA�e��ă����(���� i�ܹq'f��$]B,����k���m�sPD"
Y0�N)A�ƤaYy,�AVE��	�C.K,���z��A�b���]�ҡ��
m��~��D��V{��0��e@��j|:�YB�3�����A3��H�!t�-���!i��&��-�E�%�tCR�AlE�������T�3
����F�!�bL�������@�P۩:�&�=c4S�o�Y��J�PlYg4bc��ÄV
h�X��n�q*V���(JǴ�(�)U9�.��UASxW!�iB�Z|����c�\�U��S�l�3��u��`+$��G+*�R)ht�8�q�Uh��҄�X�ѮA�:`���^㦨f
��,TM���P��7��F'�b�SO��x%B(��T�.!֟%��2��$���~�,UhGL	*�E��+��$T�P SS}�� �]�P���@Ț2t�<�r�j4�Fմ}PM,J��;�
�j�4��H��um=�s<A�k#��3ͷ
��	�9]D�����n0��}�Bږ� �a�`T�ug0���ftu���V.cд&�(�c��r'��UqO7��&V<ns7c�S����BJTOC���U�jD\����F�&I}�����>BV�S�F�������9���Pߖ�ҥcqf-5�f�Ѵ���x�&J��(�4J�������/�5:V��q�ش�]�_mkǺ�BM�&$~�u#�_�Ӝ�[�[�Ӝ"�Ѳ��
�V�ޫ!( �x|�Zc��{m��q��B[E�m�|�ΜJ�:��;�},���j��&a-�8��p���Xo�����G��ci��iʉ$紵lh��*mg}n[h��6H��#�!lA�%��-�~/�<�H�"3ꋿ�C���A�*�3��Ec;}0N��	�����V������X�(ƧY��YBZA�*7��nz���G�z�/��G�/~O{����j��+ė���L;ЍB7�ԧ(1�Ԣ3C��{!##�*	j�*�)���I<t3K����y�9�������Ʃ��<Aߞ�K/s�%��w���{�k.���<��_\q�.�0eZlRU��M�x2�/.�Cjz�,�jJנTk�X�:×e�ĥjT3yB�"5c�d8�El-�A���(�vs�5S?���O>H��ǩ6n%O�Y;���pYr����h������n�JSn�k�q�2&�5M-�J��i�QΓZEby�!r�%���F8*\�@��`{����c,f�hFi�I0�{�^�3q������y���H,��$��+�y\q�`���]>�4l�TyeS��c��2�I�^z����
-
i4ڙ``DAch*#�Bqa�T�����0�d��|&mbe� �����2�M��Yk����J������}�NF��khZ(-����}S3<�Q���ŕ{��Ka����i�z|lQ_�uH$VQ�nsrڊs;X$�P����?�0�P��o���x9٤.'�9y�rz��u���W�?��@~�G��_��'�+?�~�Gŏ<�Ƌ�?��!��n�
L�D򖴌?%8�P�S��CH���m Q�s�5RQcѱ�K�� +�9r�4M����:u���c��U�Ʃ��g<�a�̏~=���_���Ͼ�����I�&��C��b�r(#��:X��#J��~�;5˛�j�vQ��)�W��bb�&f	�Ԅ��)#^}_��˿��|�������ч?�����y�'>�o|����o�~�w��o�nՆ�66+���2੧�Đ ��tFbaw�*	�h��[����쀭a�\pW��x�;���58k{9�j����+M�WB�=>��͔rZP�o�h��>�>^�g�܇�7P�	�lc���������l��Z�}hU�@��y��d]�e)�B1��'L�_�}���n�;����KP��$�i*2<&Z���Z���{�Z,�]�0r��ΏF%�����Űf����k���_�̟��sy֓rѡX|"V�t��q�(�kUh��5^����6��ZwWa���3�tl[Ѹ��gN�1܄�Eص�	�<��}���~ŗ�?�S<�~9x)'��Q)�s5�h��`�|�{;h��m��C�9���}���fAU
ve9���nF3Z������=��S8v�$p��m,����/Y(Ģ	���1����nU+��Ƈ2^ؽ�@*%�W�g7�|��������O����F~��ɯ�޿���i>���Z���&db�4ʅ�]ͩ.w7o�W���)TV�n�dX1\ҌGP���]�3�}4��S��37�����������w�w�>�	Fgq��}�>��9WM�{�u�EU�bE�����U��w5�?�q~�	O�ǿ�)��7?��>�����~����8����zO��籞眞�0I���qQRTQ[�$�H��}����gd�2�s�5�:T5�t�4g�4�L��h�Oq�K���=�^�{�߱q|U��\�-�"����q�p�A�>����5PbP��S箥jD頃�	��$iJ���'Wwq�e>}l�O�Z�C���˧F\w����`�X�!�K�:�#Mzz�������W9}zi�����M�f�@���|(�[�����?�=/�s���u֒��im���̴�"�d$1�L�Q��[����0�����m5��@��R���tO��3�H?�	���.>��W�7�26?�	����=���D9���B91�f�Q���s��{<�VjUh#��,}��D<6Oc�4ac����Fg��۾���_������?�~��/��^��G!�k�U�I���`m�t�2Z�Pt(r�gZ5lN+���^�`"p��񾏰D�kU�U�@�]����]�I�ڄѫ��/�/�={s����ĭG��E�c��ńG?�*.]��	������X�9@�}٬x�'�qblYw�4QI*��w������^��<l'x��rM�l�D#�x66��%��q�,����{�[~Uu��]��ۧO2�$!���@h��(��ł��������(
�PU�:��Rf&�v��rڷ���c�s��$3��^�=�;�{����^{���g}֣���\$7}�3����C���r�`I�,��d�"��-2}�gdK���V`�Ev<qS�Ck�T/C��������������'�3l�7��d��G�t|�(���X�7�H��!Lq�np0��s�L�f�^8К���}�.kرc*�����܎7C4c�(1���Q���c�p*p<4�j��Ѧ��=��=��$��u�xӺ���Fp�i�EE���vı;of��y�cw�#w�|톛5�T
\1b��b��=��4˦�ЖZ�Z�^hZ٥Nr�$����=!yҊh�HC�<d	:���'\eXH��jO3eA�p�G$�1�mG��X��:��sOɖ3@��B�S"�	Cs����N<U]�_[&ݴ�s��⧾�>�ѯC����
v�g\�E���l��mbR�,ų�O6�a<,�5$B08q�v"Ie�5.�k$�Is�d�=�{�==D�U��|�h��L�F"\w�M���"�2(�#^� ���9x�Nf�;�ϴ�/���;����7�.Pr�{��&o���n������m;�
����ن�tB�`*��wJ�4��7��Yȯa�,k�����/>�5����ͥ��zs�6$+R'�V��H�is3S���9����x�ԗփ�)��� ��RW��SG������p��g�T�EV����~S��~�]8}.�s>����5eQ��"�@kA�*���GHY��(l��� �o�N'^:_b�@�d�$h�OPN�x��e:̷�����~��W��+��~���?/���mtV��X�*rp?^��+|�U�8Ϭ��[֭�{�}v~a��{|:9v�����"k�Gy��ϯ~�s+��l�_�ߗ�+?�8�����͏2�Q]w�9��% Q�� PǾː{��c\����uy�8*=M8�|��|����c-EUb�#k�B��ш=��+�v�_��D�սY���x���A�;��+W<�Kz$cK���y���*?N+:0'N���>��C��M�H��{��%���X%H[:|@0����&�����/�Ox�E\�O0������8x�$��b\@�ը�U�V�Q�c��U�f�Ŗۄ�p��)6��cD/���To��IB'Kɒ�������w�YZmX^�w�EO����y<��m��Q���u,	�aM#L�z�ڣ�!>쒠#�҂�@��+|�>ʺ!Mr�Ds�9ۑ���/���|�o��<���~�9����}/~�#i��?L=!�I��Е�,�4�Q�|���q�$I�YJ�49���05��x ������1��ů��_�2?���c�c.�S��{����p�SR�mf.����KQ�~�)[��-)7�H"N���-� �gY>M5�V��r�z��V�g=��=�ȿ�3W}�����۱4T!�A=24c�ơD�С~�3��w��4�f[��L��M�x01��J��4È����s��/�{�������_�m�x#����s������}��x�B5�X;��5�0a�F����4�d�L ��AP#E�h7�R�!4uQ3�m�j��k��/�	��O}z�_��z�����y.�O����~	fm�z8ƻoKT=��j��M ��l�FM�.�0��a1��4�DK�CUB�	$�EB�ړM��ٿ�~է���^(�LP�©���)�RA��H�eB@�!GL�|z�hl8���l'�\=��^�c<`�~����}:-��%�ՃH5��xs3��x���[1v�NW��)�C�Rt�P7g7 �iŞ�p�*�D8�Wc0�V�dj�M�O~���m���n���$��
���5��[��+��y�r_�w=�!`8Sb������F?!.P��9}��X���%�V���Y�gP����+���+y�?��������(_�R��~�a�LLEa��c�8g�A�{.��TqqhJ*Ԣ(PJ1??��0q�g��K�p~�!�e�_Ϋ����G���߸��O�=�}����s�p`u�z���@eYX�������ϑg+�ƪ͛�_���ޣ��-�^���]�9�X����{x���c�y���\��HU8��ޞpك�rߋzt�>�r�E+p�pH�L%V&Ay�vAL��2�a)<�|�/�/Ρl��{ ��r�ލ�y W]��}��
�H3�������\�('8�A�(�B�,ڻg.n]�edaI ֧��aYI�.�"I`�����~hL{�b�^�8\{?���!��c�EYöi���$�cl�T)�Y��A����k���L@	�&�U���j��r����Ƭ'�W���gk.5kj��~��� ������h�?��x�X�0�K�,E��Y`�����B1����Bl`N���48w��g?����m)������7��_x�S��_~&�{��|:3�b銇/�ۯ}��p��eue���ۘ�
�!i��-8� ob��z�]!Q�uV���Ga;81Gm{�q�����t����mq�羶L�Z l(X3I�L<�Z5����!���i��X��FH�����(��
���NiR:3{i�Sa�<�\A�P��{�L�PaLjJ�R��<���aﮈMX�d0����J�JQ��e̶ڴ������n���r��4Û��O|6��s�W����
�GjMS�u|���l���Y�Y�P!ˇ\G)�铨����r@'K�5��)��{�9�L�ޙ��:%¤H����f[��:h9�5=�� �A���BB���IϠ��H�H�n-<-�����dJ�����s�K��i /;Q4X@(=���y#C~��	�g%���~C�p��2�g���Xff{h-9|��u����N��4>o�6lpt��vFuFHP�%�8�2n$FiT��ҳ_bN'�n�C���4Kq4�SU55P	��h�x<f�3Cb5�KL�*aǹ��i��/=����ξ����J�T� "�g����9yE�I�Ĩ>.��>:W��3a
"<�t:��mv�s!���x��^�O������K�J^�;��/��C�����[��*V�<	�/|�W��o��7|�k�~���]�ζ#+�CJ��2��3A&߻�р�c���[��+@��NfW�qi8̈ft3^BTKL'�-K"
n�拴Ԉjt���G=j�T�@�"�1`RƋ�b'q^/"h"�c���*�W�a��# ��""ċ�Y�m
��`�?`i�@��q�ۻ��`o*z�a��w�zx	���Ɠ����!�<�s�4�H��|Nώ�A6���_�OX�d����l���G�4�fU��K�Ul�":J�2 �=j!YZ]�2�i�0��T��`�PUϚ ���`^�y�{��1���������՘�l���{)�(4�+B�b�Ж<�$�g��V�	�(t���qP��x8�hI�ݬ�ȶ�u��GoL�nt!W~������|�@������w|�ִ`��������7*��@��e��d�7h�M�Q��(�uT���1���H�9��!!�դ&E���e�f��H�S��-��2;��f��D������$�c�of�̘�<h��4��2i��_M�4]YK��l1�Y�Exݨ
˿F��RD$�R.E���:]*�B�0���Q�������4�Ix�/�V���Zc�tMq+��{�a��/��KG��3�yZ$�(f���q�B�AJ���x"S�|�}x*�_`UM�@#Ά{��d@9\c�ݣ��2��wA�T�1���0�-VT��x�������54}��O�@&<�$����D�w���F���>�07I���RA����Uk� blУ�P��[�U��-t"�}���;�i�w"�=�a��J�#���s�J	��R���nF�|��>��\��� @쿽蹋hm��%4�����4b'V���	�v�ɹ09'Ρ��y�21e�)�Pb�"�����^�^��R"Eư?d������/�/�q�~q��=��6.��x��/�%?�l��O��O�ĨR�!�ޣ�Uq1��v�=���2��N� ��.�űl�R��4A��D�h�cj�Nn�s����4<���<�����9�%37s��ws�e�����UXƦ�	H�'�!�(��H��3_@y�h�LDDV԰�Ŀ���*lB���A#��G�(+ �۷��g\ߔ|���{;γy����p(�,~�p|�)ȥ �SS����#2%	�uc7�װ�vA�ʂu�yȖ
*�p�`���"l��qÊl6D�X�bD�Y�^��s�!Őrk�݁��H{���huqy��2�w?�.�c��R5�T�e�
�/-��ZK�V�\Ef-ڛ`"�NL���܉�h��L��P&�*ih��L�a�Q~3lq�1�o;B.������S���o~��G��_�t������ǿ
���s�J�K��t'��H���KPF�9O�2W���j�w訨�O�i��V�'�bُ"���	����6D���̰RI����� k�k_�^��G�߇�zѥ�苮��R|�(���_b��5��M&�X�0��0ED��@�5!��^F�!k���S�@f%�IR��N��$�٠"qΰ����7N��Ds��>�?��K���-���k���~��}�o��Y�<�W_�G��v8p�iki���vL����1}R��Hs��9p��t��P��I>���ʖ

a9IP�r �O�D����ΆA��z��a��o�9�c�D��2t���9*i��{�l
�N�9>�e�ǿ7�6��.2����r�C	�5��(oP.����zJL��sB�� B�&�| A�f�X��Е%a��}�y>��������PJSG��p�Qxǿ,�W^ŗn\���^�d�3d�sx�Z]8�(o��� �Xe���dI����_x��al2��2������-5��--��B&�Ɩ{/a�Ly�{?��7��u!?����=Oy ۶�ܲ�� ����)�4�e:�Y�H[��	�u}���7H���B�@&B.�߄�&ζu'2�<���ޢSE�h�u�\4;�CG�B�4(3����x�u|���W=�(����B1���4�x��X�sI$'ې`�D%�tn��E�i����eK�Z z'�0��LtS�69-��$5
�"T�b]��]d��(�։�S-�$�M�-0(s��_>�_��?���c��{oR���@9�2e�M�����C�C��:�	+"�s	�� �\4έ����c�m0���h�H@�9��fv;��m�7��x��?�^�Q^�'7�s��5^�����y=����6��L��˷aT+(��$ޢm�r���Zj*��TB%3*�P06L�x��C�=�{H�]0�SY:$6о���P@���T�����>��[��w~�w��O|n:_���}w�G�>�_G0�K��ٝA&)H���R�SH4�4�o�*��sV$���FOL`t5����,VY��Z--�l(uC!c׀vt%��>p����u��Ӿ��?����c��۟���O⍗=�������S����\�d_m87�*��� ��U�0@Q*A���:Rv�'�jD˟ND�)�x������d	Ѵ��^X�6�1�?Yi6�8�C�j��^m��
�}�A	�����Q�|:Ű�ptM�<��:�4!Q�/r����g	U����B��ͼS�9���+&r`����S����hw�b@�{�E{�b�����N��v)�+�_;Xp���S{h�����"Tdg+,^9��a�JA-�T�2���j�ݏ�O�'��NL`1�zƝh���p��	�¢uF�H��n��{07����2�����I��>��?v+_�FE�β�KH�=�4	���~���$��|=�2�T�&si��2�d^��#�s4��
��P&*��{oi'�]�w�ȏ�}��3s����ބ��&z�����M͞��|!���������⼀4��������W�%�	��^�x��L�ߎ��t�;3��S���
FW�DO��b�~�&�tB����ę86\�N���u[�X�&�jg�6�.a�Ye��t�.�1�+�h�4��31��ā�a��EeY'����:%19�I�F�Z�\C�K2W�45��^2�lv.i���*��i�{�ڹ���YR��<%u^Ҡ)EB!J%��ѡr�aBSX�#,<���P ,$��(�Ė����|8��'Y
J������k���h�����;�a��MKm��|z��Mo~�V�TV$nxr���&8k�cm�r��"���8��A6q�+��*���G��5-�(RK��
��+̥�#���cv��v�Z�)�|U���р�(S��&Ĳ�%�c+p��v��dZ��]KZF���mz+�)�UH�M�J�W�3�-T��c�	09��Ȇ�;�{"�+����M�	q�4������V�;�[�x��
�-Mck�eu�p"�ݝuP"A�fo����@H=9`�>8��gԀ!'���q��x���-�N"�G��l�Y`��W��3ݝee�$�͓O�@���|�6-r��1�����[Y�C�'#��z�5X�N�Dl��nǣ�ug	 #7���7?p�x<�����15�V(�Q6�����l#_�Gkۅd��q���E]	r-�U��Khl8�Nΐ�bmC��X�X%�����o�T��֫��!|0�/H�$q�� M��T
4��5�񘶃^%�=Y��SY�f6UL%g+��(<-���2%�q�#�b�T>�>!�,��҆>���#���zmUA�G	������>�[)2	[z����#�WY�%������,ѤZ��D���)IK
Z�c+�"�6���N2��U�Lj
+��c��I�V���L���"��n���N(��!� L�R0=�I�b\9�#(��e]lڡIR
C��[/QI��(��oٶ��<O�T�Le̴��R�5)=7MZ�l���P�A*$J��֒D+R)b2A7��f��-/����v��%�6c�,����[]��B��Ti�[	B��:��И�N�83��"�n'����{CiƠZ�l�Ʀ(�&�)��1�S�.AxEc�tP�$�ftڊj�J7�R�r%�S9�7�� �@;h)ȥ��3Z*�z�cKb$�x�� Zdx�I��F� ��ř���֑��Yz�딮ɘ�E�Q��46P�����d�h���)B1�CACI�Ԃ�)I�l�N���4H��z�u�rw39����$��~�M�l���?�NFY���jJG;z/��NG�wPD��$"K�P�-�Y���*���7x[��C�ki,X#���T嘪1.��Ǝq��a\�\�!.�d/y����o��i�07��zH�R�&bPݙid+d��u��5(�ΡՅ�4���.*(J��Q�0�jFU͠)�c�14��i�n�i�j�6���X���ፃ��k�j���n���O0�isήyF�5�&(���xGk����~Q�w�h2Ih���F?����t�<W� k�q�z6X�3�6�T�sX����5B%붥�	�L�2C�!S��>X���Ʋ�2`�ۣ�j�q����*�Q��x�V�T�GJIa�0WLø,�Ra�����V22:�it0���E�(I(�V�r�\0ŝ��i���U�"u�r�L� �T�!S���H�����s4��KG�g�j7�-�{�D�h��:�*��=W����ge	�>tk,diK]9ʢ��B+k��
�$']�N�:A%�4l	y*I�p^J2I��״�u���L�P��b��s8t�qt��%�^Dgv���Y)�F(Fe���GC�!)�Z#q#t3@�+�����L�����<2�jD����pY���!�%p-0m��P�un�y�AIK*�|�4�M�.G���ݢ_@�3��9��~c=���P
�sx')���Ga*�t��TF���LOo#m��+ϱ�1˃��
�O�>Ë)S�H�B����� Jl������J�0ģ�4��b�9u-i�4�gJf��MO��Z�s�r*��4:����6��Dw3���d�Ya�r�� ��$d�~�TKr��saIi��(]AZ����C'j���k�O2�n�j�d-Z$��W�Jzl")�g����\�A�JMOu���'o)�����{B�T�P�r�1;�M�B<�+���e�:h�s8o�f���B�)J�$d�i�H�����+�+���|��M3��G4� �܌h�
S�ت��%�
�j��a��;�0�<����c�7^_��˨z3	'V��q""���.Sݜ^K�o%W%��:%�����2��
U��3#��l��%�V[�*f�Ę!��i��(����5���CQ�7S�h�>U=�?s��א&`�>�h��nF90C�;yS6���5�n�T���1$c�+'8~l	g+���Ne�#ʺ�i��\�Z*Sb�_��z�k�8��[�����M]��]���C��@���q�e�BY�Q7#���2$Y�gUM#ai���5�X��tn�2S�N�g�%��2����hښs�z˚0���eQ��cH8�T���vϪq�Ǫ�XǊw�:�H(V��Z4IB�y�q`m��5�b�"������&�$�p�f}9C�RA'F�!-��uH��4��ʀ��z]��2���s�I
l�HS��C��8�.�?�`��5Ǳ&4߄f���f��Z�TCL5Ė}\l�X���0Lp;��!ޮ���b�5n��Zp�Nr=`~Ƴs[J����9C�U��Z���d��]���q��;���!�R!���W����:���	d��*V��*�8�.�P�4'�	�YB4'P����I3F7c��X���,2=Us�gP~	Q�-+w�m*eG>�����&	:��4��:x$eŉ��c�U����L}��`�J���
�����ތ�v�w��؂̖��O�����[%sCW�ʆK�4������=�Q�UW�eC58�Tf�iA;)�bm�V�Ԡ�(�'H>�|�3�y��`n_qx\�w�2I1i��x|ҡ"��9���~��D��D�s��s���H�ñv��<g-O��FfX٢-*�b�3�i�j�r"�,e��b�v1�4����nC�ncU������i���gi��<Z85 �$���Dluh]ZZz��ݻ?m�S��`0�w��|�曑^��+��?���Crvn���;��?�~����1������Ӂ,�$�Ň,~!H�l}-�pz�UG�I-R� ��e�r�vb�JXe��`)�H�8,�S���m��\�x�C��c�w�|��x��01;?K��Z.��}y�G>���Y~�7�ϝ��Q�H[�d�Y����ok�7�~_��f��M�XRo��v���F!}��)B(�2���p�S��k�n��v��}���}��3O��
���πH�[]�����㪏��ޗ��_� �W�R��6��a\Z��Yfg�)FE�eMadL��-H�D`��	��j�qL/�0�+���U�c��b8죵�(���h� W<�^�򥏥Sz��Gp�W����y�5O���׿�K�>�i���ex����+�D3�J�Y۸u�b+�V!�`��
�� ��e,��!A)��4��S@lMԅ!��jk��bٖ�����������'����U��G��j,Y�0�$����_w� ���j���'�i�t
��]��\e�WB�b1��]x.��|����J���/��J)F!���p�\ʟ��C�{�n-��{B >VZ�1;~2���P�f� ���Z�@{��Ć��Q0NBv�����ѡ,�:���b���-�OA3X��;��c}��,L��k�h4�t�������4,��r�MX/�z��u L��N���un.	ica�Ф�`�耋1X�A,�+f�3���=�3�N��.���_������9�KF��񵡶%/���W��;w���/\�t����=��͉����l�ߎ�.@�	%3�G$)ބ���Ӕ6���5N@EXR;)��`��H��4AUY*S��y��;�s��a�*x�#/���}AB����c\ig^��W�+��J8�Lq�M��U�)h�sjgq2�Ǥ�tI��P�ر�٣m����%6K�T���=�����P�V������5�aREr�>ر�׼�w��7�%d�O�I�r��ӄ�큃�
���x��]{�r���.8�[n����+��<���	�8ܔ�^�aY�ޱ��������αY)���M��}�$�h�o�8�	� �r/�7�6O�ƣ��@�����0?�}�
{����,?F����R�C[sޅ��K_�**j6IR���Ŝ��!@L��5H�!!� ��M''(���L����&�z��<�9��X���/2��2X�92���)k��_t/���J�~J����@����3B	����a�m�f%!]LFa��0��o���4�$a��%a��q�|�O1�)�l3(�4x�gfY[]c��e��s��?�����T3�HFD$�F���**�`ʎ��E��XNVM�.�sD�Q�UD�Ҳv��?�;���%���9�T���-�
�D��(�����k��O9G�y
A�}�]�7n�\��w��|P ĉIZV�i���ᶀI� ;��t1�d�P�l_���<�R��D(��b a#c�B����b6H��B�' q6���
8������?^c�L&{Ԟ͟��B�c.��M�����!ȀbB0�N4X!i���K����Й����Y]�#�N�ا��P*�M2M&�ǿ����J�'�4����2��=v�o���n]A�'�Xߙ����YGHm���ub��=�9>���s�{7���)�#�N��\��JTT��jC�uX  �����������ȝ�v��sN�����?�bn����+�������[�E,[�!|�F}���x���u2�!���s\�@P�bE�/���5aNz�>�6�Y�E|ZQ6����U���@c�^�H¢�"}��^�4(o�r�u/���$�9CS<-i�RV%lc�	ߓ��`���C��\E"�	,L�RtH˒�#\�I[�R�F��9Nc��c�L��O�v�}w���9���P�P\�֫���D`jO��~��AQ���g������Y��>i��'�m�� �i6Ĭ
�C�*�w�)O4]X��^=��f����Q�p���z���/1R�'~�bOm3����M����uW���It0m*ի/��#�> ��8
�&-������>��j�ST� ʓ���
��q�`j��dB��GP��H���N�v�s�������7�哣�#X��6����	���FF�(T"$2x�:���?9���2��*7/��pk6d�lŰw �~��͋Iz}D!�ͫD�P!r2����*4r'ׇ�i\^�^��{�_�5��	������X��4��vW!�?�%�)���C.���؊MY#��MU�3���V;!˓���7���ģ�	�-�I"Щ��$)ZX4�JɅ>kF1�%�X~B�51Qb�����ucʝ��&'<F�X�)��tW���tW�͇��H�~*Y�g������n�ʖ
�2L2b�x��h]&&��.���y8��g�l,� &H��� ����.7cD��M�F��≩w6dH�^W���m~O ����7���4&�)MȮ�-�2Q�}�,Jid�ij�x\3.jC�&R�&�B�6���8�q���1ҷյi,i��j�Pچ����JK�OBn�ϱ"R����:x���=:�@T:i]�����ܛ(8�D�ꡣ�L��E�Q�w����NAٜ��6��𓳀YA97n�	|�6��w��m�����vw�އ���t�Ý�6��$�'(��a�&�Q�N�I1�����S�Nӿow��G3W�92jL4�,,��q��-��$%Q)�pT	���Z��Y��k=�l4&m݁u&WЩB�I�2#i��#���@d�5XMx@��.���v��E�X*[5�d����".���9Y,<��b:�!@1y�Y����G┷8�I;h�q�Z���=1!�7��O{u���@����-�C2Q�L��fRH��\J�2R�&q9�OIb�2=�<3!I�4ML<�'�?,g�<�D��xzx�!�F:��
��8��D`c��OqT�1��Ρ$h4�y���P��䔦Ш�:�yq�[W`8P5V(�ʱ2���fl�!=V��i8�N���a��ɼ
�d}��𛬒���Ǫ��z����
�n�����'���~����N�����wx�	�Lq�ܬ�~����l�yګxyfW'�V�Z
�p*�-���I1,0*'�$n6�:�Qn6o���mr��gp�!{�T�uB#5	��]�c�lJ�j2�-�J#�����8�Sn��ÞR���6�'��nP�~���(B�����r�&�sH�ud>����<d.�X�B�=��ޓ{O����m�$m[��:�ma��ݎ֗ L��y�a�޳�e��رc�ܳ�OY'� |�������[�x�����B���p�V���cT׈��c��8��ַb}�ӳ��m�*�@�NდE���(����ԫw���ciu�=��E� ����������w�_Z���n���d��.��ǋ�
(�{��������t8�xg!o�����(��v�cqA[������g��}��7Je�L�p��ؿ�.ڳ�������&ue��`4�¹���ٵ��G������<�
��=�qU���=�Q��c��.��̉��t���v�{Ϲ7k�#�;�~��|�s��^�h!�fkZ��x�N���!�0O%�x����g=����1���N�CQ�!��Yb�sIB�f���@�����\�(jfg�q�&m�����⻟�lFu�9�S���X<ZKZY���2B��=@�����v���_U.����
�DP�=���R1���V)�av�n��������'r���llL�_��]f�)��Se���������0?�(��(�o~T@S��2������<�Q��O]��!	���3T���,$y�d]�,�%�	�&���ȷ꿕����@�@j`�Π/����_���IB�{8+0uCQ��Jr�=�O~������;(~�����"} �p�$,0[���
�Q�7�~hY��<����}��"���֚��\������p�8�M�4ƅ��TK�	z;0y�ayF"7�:�tr0U�
��~��^�_��m�&�g�J�$������Ǐ��=�\e�W�IAwq�7n>IA�k��ʦ�v�W�����o��k���G)��U��&S���*^�]dr������״�yަ�@����cx�9�'�k�g�E��03����%fv��k���)^��O�#5u]3=;��	em�R�fUY�O� h<��L���10�1-�9o�~t����S�]��q ){Egj��p�^�"^���E�M�ώ�馛E�r��f�����)��`T�`�UN�'_U�&=�����t�17���o?JQh��m��} �x���s��_����"�@<����� �����i���?���|�i�3�n��:(�HU�A�F? �WH��3���Ph��x%8Q�Yi*�����?�rVf�<��~��^�Eڝ�q�S�<O��{ ����.--=|�6�)�G��-���=\����2��W�#?�#?�i*\3 K\���k~������\�rv�s�Lr���|�rB�?bb�?���UxI�Z�g�^�q����3���|(Oz�4�)2o�Fq�&�W�������w��߿��4�V�V����h���ũ�ޤ���6�w�
�Ѱd׶�Hk9|�7�Ϲ;X;�ut�W��I���oᵯ|��I�P���,�����^����?���C5�;:�H�RhVW��v'�)6&rTTO0ѿ�&�-C����
���HrZ�"#~�*y�9��?@=�\���I�Jz�F�/�ٗ�[��|�'����$�3�椵#SV�iJ��F ����·���ҕ\p�ZR65U&9�4��4�<�;x~�7���˿�ZҴͨ�AJv,p��R��ZA��� �;iU�;�z���!I��R"�"m�hw�7�;
ѣ3Tr�Z͝�*9�-[-f��!���Ջ)�m;�my	ѝbjǹԲM%R^d�`���XG�O!ul�w~��p�׮[�_�9�ӳ�'�Ցbm�Y�
�ٲU�y1�M���W�3�/di��8JIz���7N ;������x��^�PL��ڪb~a'}ĥ\�����[�`v?U{7U{/E��Q���w�tgl��;BKB%ۨ�v̷h�X8m��v���rV�U�<��9��{s����j�v�Ci%hA];�׆t��x��?���zP��5�t�h-s�f�f�fJ�L)����ϳ�d���������T���N騊���K;ښ{m�G���C�y7T#��Ǡ��ir9
7*I��dY���VA�_wݮKpl�ZO]W�D2�J�����>,���N��Z'�v"����>��'�������ZD[_�h!dk�+2�J��r�w/0�<ñ�՚��h	{���U5e9bvv�������]�ϣ�[ ͦ@��[St��!dC���ΦNےt
�c8��{���:�1�λd;s��a�6�*�./.1 �IZ�$��p�׎�VBE��f�LJ�[*M����R�VljZ��i|��wU)�*e\n}j��W���}�O�cC�2�9U2Kk���.ⶃk������Y�H��,�)� mf��YVt]�h[ G#Zΐ�-���2Ӑ��n_SS�7y]����7�a���-K��p���>����di�B���#7���FN��A���B@Ģn�I�L��2�^Й���,:��j�i�-:�.�M����3ZYN���>�ɓZ�i�L��[_��"��7][�5�ݷ�#��ԕ����			p�m��k�6Rk�GA�9z�V�����4E�z��N�C�$�z	��4E"J)�Vg�����b̽�%Y���k�6I�033�p�;��H�h��X+K����\w��j���\d�2#9�$���-�CK[t�����t���S3[_�3����+��U:��_���fTF�LJ;�c*����јV��#|�+���ѩE%��x!k�@�
��rC5J�&e�RTH�UcP¢�w��a���B"隊)W�iD�i)�3;Ř�K��%��T�����|�eKu�	�\�x��&�$���<���x`����x �k�P��:�Lj���@�ļ<c�U��ԱU~�5���ui0eMU�TuM_ך�r4��.M�(��u�D�ꉊ4͙��b�?�IŶm��z�i�����)f�����U�ʐ&9������`�w��=��0M��65S7��������C��є��]TP�0�a�8��QU5���O|�Z<��;���c�����ׁţ' Hu�R��'X҇�B�J�L+�$��D����4�qk-u�i*OU[��n�z�ړ$	I��O��:!M���,.'�2fg� �Z$�)�����Y�`kC"S��R�e)�v�o�W��H	�na}�'\�N��	<25��Od���T�+S*��[-����1�gdB"M��К�1(�I[9�m�]�܎mT&��V�TP�}(��h����FFjK�J���U�v	t;m�m����������/H�en:A��]�V%s��CūTI�SM�=u5$Q�v�ޑhO�x�hՉ��^B����V+eT��ٜ�fD]�0o��4Bj|�鯎����Q�����<s=E�Ԩ�D�'��|��d�#�<�b���^ȱ�N,�v���4��\3���D0�l>�S��|�s�9�B8�s���*��6�\�tw���6��}�0�!&Q�5��`��$�J0JJj�K��h�PU^+\��T���q's��j�1XSQ7E3��ǘ�D�����49-F���qX*��D:�Qէ����	��5��XM��ƴtE�^�li\P���iT`0"���y��I��0"���ӌ�,#�t506P��{�Z&4�l��%���@���F�<^���G�"06���a+C1źC���E�g)[*����HDx B�]k��m��¿��&��I�/�~ʾگ@8�����Ո�cC�oH$4՘�h���<S4���x��5�&LD���#%Ș(/ ��'\��j�#`�$�`��qC��]J����u$JGDA�X��rL�_��0\[��)��x�p4�,kc ��n�fېx�U��&d���ķJ��,�S�2� J��p�a#,Q��t`v:!MS�����+,M��{i@&I��-�JQ"0��h�vH�w^��(൉)d�N�	8qD��l�
�F9���&�H���<��QJ��2��wHӜ�xL�7�NZ��E�����$)+�s�3RО��3�Ee	����uo�V�nA�d����%,�c[��\�'��-�+��]�}���H�eb]-%*O!��L�I3�-��b��Y^����S3fl��Ոb��r��4H�)���XI�������������Ê�F�������%h2�l�T�L���d� �2?b6�Q�e8^�f��fv{�'�NנJ��I�!���zTH�9k	Ū´r�cԤ�I �RΠL�0%�*T���Kڀ+�d���ԸjiKR%I�!'/�B�"H�@!�(J�(e ���8Ѝ$�	I��uN�$��h�cL�m�8oh���;���P�5s�y�Ř����wچ#����(Ɣ"���G�4��Omk��`����A��k��-T����g*bc?�iXn��(�	O�L�JK���c��v^���ϱ=_ᜩ1��������A����8��E�w���wx[aMqV
���}(�G��> ӵY��Ȑ#$.�\;�|6Ƭ�Ĵ<�tzio�\�⑫YY�Y��"��¢�d��ݔ'yV�Bv!}.���y^�*��`T,R6}�\�%��	��8��ts�9��ퟥ�����-�F$i`R���D`�1���M�Ӊ��^��ً���}�w�*���(˚�(��[��`����t���Q,���FSr�k8�kqS"�J�pm�p��qU�#ڭ`�HI�"@�ZN��
v~�cR�o#s�	�c��0�:H3��+:��u	�~�.^��}<�I�������X�ُ�ᇟ���}�����=��x������C��hJ	�y�����w�ġ|�u0��Y��W���4Uh��'ne{��/��W?�����x��<�W�̣y��m��4+_g&�q�bl��g+� �ĭb	�3����O2�bMK�NI�I�
�<õ�T�ٞ.r�R}?����<�~�^(���,߄#J,�Z$X��Ry��m�Y�@�G(�FT�<��1��v���`�X*�/:��������/�^��?���!^������G��4�ޗ���V7,�+4-�b6M�ޝ:��������F�|���u��1Y�P��W����k�����y���sx�3/�i��牗���'�������<e�g=���<qOz�N��J`-�J�:��Lir��PK�O�Ɏ09�j�9k�Ŏ�p��gx�S/�E�>��T@��A{�%Ϻ//}�cx��i��7#�1��"d_Ee�"���fr�z���&�:U.Pd�,K����z�ұ���;�t��<�a����Ͼ�2^��G�k/�N~���{_�>K���k�4Ά:1~�aC���EB!=���&6zk'���.��r�9{0N45�L���au�?��7���=�~���<���}'�n#{�C�������x�^@����	Z���n�Ƨ��D���ι-!�wW\4g�)�q2�e2�����3W��"נ�u	�
�X*��%á;VH$)|��F%8����#ɶ�i�bvC4�d���br�D����0-R�s����x�m��O}���U��oo��^c�C���s}z�c��Y5`�pX�P�5㴡L��L�hb�j�EyH� 3�����d�$�KY^0��ҋ�y��̓��,�a���g<��{x��/f�'-V�uj�%���[��(��Ǒ3�{can]���������}�skQpK*����Wڏz(�w4��/|�O�������S��\� �P54U�q�A��V	����g�S�l�1qu�ω��u��O�I���n�����^����o�8�����y/?����ӯ�+~�g~��~�+�����܏��ꆳC��TpJYkijKY�E&æ���:QN)l������4��Tr�p�ws��5�����Y��������$���/�w�!��ݟG9x�#��G=o�y*�^E��7�x=���}|��T�d�.�L(JC1�0��؋y��������?���Џ�?��o�s�]c�4<��;��ҽd��)pnR�:XK2>�Fz�
�!�����y�I'ey8f۾�|��7(fg�������_}�{x�3�ū��"�����?o������4>��������왝��4�	�,��P���ʖ
���%wA��v��y�R*��ܳ�A�#�����36]���geq�p'�}8./aԺ�G�]�`���}!}GGp���e�J��I��(s)pZ#�tB_vڴ*s��8kA�s8*t�N�X��iť�Đ�#��� ��h'�s�ϒx�)x�߽�O3��"|g_�����M�Xk8��VN��1*�q	�ָ:E��v����ocL�Z�

���Y2��<Ι�MtֲV5�4�Y��B�Gx�ePy��U���}۾�|�CX���?{K+0׃���!�E0$�iPIX	��,I׏����W���aa6�w Rذ z�u��q��;��qM{z�k�/~�~λ �67����_�o�;�w������g��y+'�s��nd�U��*���Z�R�!-�[,�I�����x<i���	�R����2��i;��- H�D�F�P�mz�d#��cŶ����pߋ��\�,����:5G�r��,� �0�g(v�O�>Ax��IO�U=�qmx������i���$ֆ�{�.n;p+���[��3�e�*9�������S�
��Xk3�!֩��\���O�WU�����롬J2ӹ�O|xH�����������d'����߼�*�c8g/���#�ƛ1�:��|`�Ф�0s�#u.����'z���!91!{=����}��ۡ?��o�c�%γ�����uͽ��{�[���8���ܔ(S!|�B�z8��l��K2����d��q� �/���sHoC|��@�"T���V����S��4�)q�~໿�^*_�ʍԵB�%���!_KE��م�%N����X�^ \`��Bsby��w� �1����u�.<��W�s^�z�:���=�s.{��1'�p��C(�'a��52� e��R`C	�3��9�eQ)�"ċe0};�LAj���σￇ�����_�a��f��w��6�����k�[�F�y���d��$h
��Ix{vGtjG�1�vC1' �j�VUT�f�^�����u�(��wp�v��<�À�U��@|WB+�����D��$���f�=%[*�=ݐu�K�c��(�a*'Q>(��)���"C�P�wi�({wN��e |�w0692�B���H�K�Er&��������d�;"$
w�]fff�_����������<�=��-{�*���G�����#;�g>w-J�#LѢ��	�3���Y���6�"�t������*pU�0�&I�U�ض�����ۏC��,�:��3KY�ܾs�Ǻ�C�z�3'7�Q��xH�'��������@+���$�5%�?��0Յ�5��������ۚ&��Dx�TQ��jh	EWh�2 �E�P��pq:����@�6D���.�N+I��eZV�[Aրv���6<�i��I����1z����Hd *@տX�b�	����fD|&���Lۉ㨕$غay�`�%d�S~����;�r ?���[?����Ͻ��<�"|	����}��Խ�zB- ���cc2�66�V��!�`�w###z|�tm�IuF�7�u7"O�ɾs�c��2��K7I��k�y�m�[؍�`Z��^F�*W�xNa�(����H�l$���4��E I�(���45�������r���b8FYO;k	@��(R����?k4��BQF"��i9]�Z;ב��bTX��ǆ)���'�@Ȱ�J�0%��҆�<aR�������-�A��D$$B����e�`�J1�Ù�р��uB+�c��9r��}�]�r���Y�y�����t�6�(������w]�u7܂R]=�����@5�<�
���~",.b}ĕN$�N���Z�2]�r���M軞�Ht���Ay�������Y~����P)�q.�m(��%��u OM���bEHаB�;����5�Fe��+�{�a;�R<�7d��V
���&9Y�M��pv�JQF��y���l���Nٳ��ce�\�2���*\m4��R�:��՘J�����>���y��z���㴲y�����h!'%��T*��$��zV�XX���
/�u�b8�V�Op��/�3���]��C�;�<w/�����X��~(�w�����=<�1gum[WXk����R���}[6�o)^8�����M��Μz0�5Pٌ�Q��e�'?=$���)~��E3w2]}��_��M�y����հV��$�D�LC�����?c�PjI�%F��
��`︩HBw80�:�n�KZ-�l���3�S\�ಌ�o�D`5�2�,_��Y�>�'eKB�5PA�s��>:X��W�q�a�s�b��Q�D�s5�����ҡJ��c�f���EZ�^�
�)��y�!#�������=�I�X1���J|����^J�_�s�R�gt� �/�!:�������{^�Z~�����*�����=��<ᡈ�8�^�7eHaR�A�,��Ycq^48لg��7�4G�7�A�ݙm�d
������2�,�P��3����y���?���3ۃ~��8p��.G��HZHp�֡D��������a
FC����3gXh%�`r<+z�qI��A����ť�G���Xk��-��4Y�C����5M�n�@���/B��;�.��a3ym�����g![~�z4��O7O!8�"£�[�sHg�	�@�hvxMӠ��n*�b�h��l����6<���ػ*\��[��<V�2��|
먕�Q�[/�i��B(��e6>d/,>���@Aȩ׀t���H	��H�F��%H+6�T�.�B۽i����È�;x�O?�=y�5���;>{�@n{<��y͟�o��k��.o�'\Lj��~De-���7�	��]X��$��M�!h�!@*��aI��xZ��w�Q	I�uX�JJӰc�.ƥ�����}����L ��ێY~�o���]�޷���uW�N��H�4�'4���<oa�1��Ь5!>.t,�@��q�IZ�3=�.d۸����(rΰ0ݥ�֧Ҏ�[��z�T-�X�q^`\���
ŏ
S�jwBZ�	���J�6�7��4���P7$R��]T����RN��߬�[�'���İjn���i���D�L���1��Lj����-�p�e�%�$�����3lr�ꐤ-���O"k����2r�NvU?��Nr�N٩ÏDi~c�w8�R@B	�S�E(���rr��6p�u��&г�S�vQ��0S\s�|��\/��������Ez���ֳ����Ṷ�t|H^�ͧ�g�x�065���L�/V{����K^����o�?����o� ���W9��}�i\k� �T,�X�m�4i6Ϗ8�����I��F�����/ �a��4�P�wz\��/����I��,��f-��d`=���8��i'e\Wx)H��4MI�
�����q�ɼ9U16ϧ���{�r��9����6��Ep�W!�+K9V���c��	��1�g5z�p�g'V,ik
���Z�I� �p�ɶ��bq21�B��0EB����)�nFcȴf��%\{��V}j]#z��B�����/q����Q;g@�����Z�2c�5��g�
�[x����w�.C�#�xhqT��0�N)�&��8��[�}���Wߖs�B�y򓞊��`��)�T����,�Zr���� �72�*��&�>�z0��5��ti��#��,�n�3ꇹ�r{�v���$��,J笍j
c08jWfS cq�,�w9T��(���m��>�6�� !�,x۬�Ml~G�Z+�D��ז�����Z���O�}��������'Izd�N�~mʰ�Ɲ󛖶�v�3��<��\����ZK��@�B[�,��)ZYE�z-���6�w.��`0	�f�[� N�h�x�t)�g8�!!@�t,�k�`�'i�)�F#@���⺻�ζ(�
|�p���_��jYm,�V�D�G���3ޜ��!�����d��$R0�(��do�F9W]�ԟ��+^�\����٥en--�I�;F�%#�kA�iD��Ph��&	u�Q��N�֖2���'�{�䴳�lo�rg��#|U��-���$mhw�Ֆ���,�k[�����68x��0m�F�f�v7�?8�N��.�����r�X�(,6'k�l��堠)-i�e\In?
�z�x��Ӭ�ɱ�ȡk>E�U������|�z�2�+����yHm(�4g��%D����<1�7)h[+tnh����]˶|��;���8q�g������{�9w,�{��3e��R|�p�!�G�oK�?K/nT�P�xb|�h��T6%ٱc��O���w����A�e|�k��=��MVru���rG�auz�{G���xD���̺8��RO��0����6��yFwEN��g-^�����Y;�Bb�R�d4���!u3$O-�Ν%�Ch�C�:�]�y�O{j������)a�x�\�cg��,ef8�($�T�{��{��"Ig�>�[�u.<O�#/~&��t7Oz�>�|��<�ɏ���8�������?i�YL�C"چ�i�H�=�����sK��1�;P���vҡ�NS�K�݉/q�r�[��w�f׸���|���vX�}e��:l�C��R�QD�]`s�X6g,aad�"��DI��F8=L��3^]dg��^�'��Wp�О��?�R^���3_�r.|��y�~�g��W����?<�Mo�!��d��x��L�N�V��{9�,��Ot�e�kn�=�C`���1���]�u%睿�G?�Rণ�����]:s��;]����-�v/"��3!L�Ɋ}�a�-Q�EeIBM��w�DC+��I��=���|䓷���+����e?�~�����S���<��;��7�>v���^Sd;��u.���$N;�>�~��Dx��%�(_G�B�UN�Xհ�_�XAKgdr
[T�Mx���7���/\Λ^�4~�G��~��,��/���Ak�"T>K�L�m����as����,E�Ȝ s�ԇ,��&���#E0+�z|�/�������� �~�x�K_�3���<��_öy6<桰g�>e]��T�S5h�FO��·]@����g��2(|ن)�!��Y�RF�$��Ӆn�~�!1���p���0��M͐&�r�7E�k��ش(����q\�q�('���zLm�Oس�"N�;|����=����ZF1wu���;��>����!>����s�n���cAs'C��l�\�P�WQ�|L�s�`�e~�6��q�aX8c�jL����v`�\��ޱ����o� �v�-l?��$i�L������=.�q��A�D��;�6��`��q'Bz�'���~�i�����KOy*~����S��H��C��&V>�I>��7����377�:T9w��ڪ���{�r��|Г���je��B�>oG�&��J䬢.޶qZ�����������?|×���Ctk3�YI[0�Ԑ�v��Fe	��d_��\H��ZS�5�Z�R���@���V���PU�)�<��$Na�T �J��(�~��������q^��_�E��
/����7~�w���Ow菱���2�D#�G42|�
i[��|���i�"�|:��*%��D��{��p��5����;
_aR]����Q�~�w���o�ox����_��������K���S�{=��钠�UE" O�v(C�Q�F�aL�[���v��"�_�t�ɦ���q�A!h���L�"�������"�Fc�G%����������_>�)��C�[�x��i��~��9���`���g��D#J����$Ǉ�9��qt]���:̥X�χ���y|:E�ֿ���w���H� \��!1�Nh���ٍ�������J�ɡƇ�L��7@�B��+�ٵ��]	����8D[�@��R�E��=�Z��=���f�f+�6�l�IwAk;�5O�O"x����BG�^�a7�,wŪ�((� 0������s
�Z�(%�TNi
�fe���Z�InY�p��͚�O�ُ��Gkj�n/�Up��D����p�O~�>~[��8�	�5��Swb�T�&sӓxC�n�/*�i���r��\X.,j.*-�j;���ʒ�h�� ��x8�n�}����u^�RA�j2�!D`&'Υ%�� l �=>I��4�гH�<�[P�����������yxwirLDe�]�J/J8�� 	>r�J)�
H��d;:ف ����$�d�&KR�$H��.�AS*K�+����%6�ƛ��%N:�ܛ� �EF-rl�ī�B;Eb2R����Dr3��q�fy�f�j�bg�4�]�N� F0�k<K-ֶ�w:��[����X�I�u|(G��!3����V�X�����m3Ʋ�s
��#��j�H˴�t��e��<�ʞxK�h���¤ߓg���'�|�����d�	^8��\��k�Ѡ�@�xe ��\
RK�J2Y�+�7�Ǩ��Q���Mc�{c���\H�)��� ����	 �_�'9Z��N��t%3�LP�զ���@:�r
郧;�cm��;�D9��n=��k�)F$xd$�N/e%�(D��E�MC*!M$Ze�:Ȥ�̦�y�g�T�l����񙊀{���@� )�ҧ����L���x\D���Ԇ3��Ѱ1��[TݐK��k�M��
��!�!�QE�"��5އ|P��'�ь%��S��.�)�uO�����u�E`5�F:���G҄JT~���++Ljq�w��ӡ ���I�/B����OX6����m��s:qj��ŝ,����Bz�J'�\G��R@.�侃���pJ`e8��A�2"$θP�FYKZK�F�O����&cXF�1mzf�{�K�{������1�D9Ib,�T$� yf��yG�,ڇ]6��,5�3G�-�x��)��/=RF�Ri��e�}���x�70���",�x������gH��ƓO�<�
R�^�,�ТAS�������^�Ey��M;�Vr�G���t
z�����PS���o.��������9��a�	����>��CwgE�u!�����cr���Jꅣ%�(ip'p6,�XDx���0S�]�u5�{�k}x�O1��9V$�L�M^ �a��|�tq�ͪ-4����8C���Q
y���A�i�@�a5���8K�V�(�$#�%	�T�0=��<�6yT�	o%X�"a�ƽ�|�+�E0]��(#����X��4������8�ф���p����A#,�;��TݞX&�ܶ���,���&���	��0�`Dh��K��X�N!�D4	4��iL(K�`�����Hl#�6�yTx�`	d��I���2ރ��&���wjoO',5#jQ`��ir���Bx�`�x3���T_Q�1�����	��P��9��
�8j���AaN}[���㺂b��F�i-2.bA�`�=C	#�)E�
R�>cDF%Z�r��8�0�a���4u�J�ml�����q��i*�h~�Er�"�e�g��@��s�BP)I�d���R	J�qX��~�K��R��Z��������G+C�ۉM�S���&���z�OR�I&eb�6�����x�K铰�rC���mG(7͏Q�D�E҉l�45ږ(W��aG;D��F�c�����$n��E�7F��!ڍ�(W"���4k��D�?�'��5$�B��FH_D�3�v��h
R_�!�i�(;@��J�ѢD+�_����vE�M��(��US����Uh�'qCR;F�2�O��F�v`�`oW��1�-H\��BA/
�S�!��<\�#4Op��G��S��VH�IФR�*��o0o,��`j�m�A�a+pE��I��̭��!Id�pʸC��!�Q�%�"I�tJ�S�:��	�$a�$�t�X+
�PꄱN(U�H
�x��F*�����*$�W
*�VT�RK�Z1HFI�(~�X����RQ{<�C��ql֕��-Թ�c!dT�S�� K;,�ok����ؑE����>όZ���t�v�F�:A�Y�����~�Q�O"���*�Jϭҵ���!�ɀ^�B/[�����!]Q��B�e:,�K�b�\������!:r��\ƕ�q��O�{���O 
�����
��Ԃ�~�[�&�N�=i�9�:�+o�\�c��� .��������蹂�UR�B��i���0=w'S�8Sb��t�t^��
�9�n��w�����E�*��[�� ��tU�����؍<�A�bFç>�~��%
��h�'��'<d/����א~k���G�.��r�GU'�"�X����Xh������(�1�!����
~4��3D�5�;��+�f�n���ڬ1����ALu�<]%���]��|��7K6���H���㙞���x/L�d�~��h�r�`�եޱ����:g�=�Z�f�5i]i�A�f%ﲒ��m�V�Q�G��e��Z�ˠ�e�n�o%�ۊ~[��k�y�(k��;M3
͑�M~����Mサ�����Nʟ������eO�ӻG��ә�Ǐ�|׮]���Kd�p�ٷ?7�|3��+��.^��a�azz���ϳ�E����/���������I&����$	����NL�����:���tER���W��k�#��g=�~L7�?������Щ�&:�P�+��s_���fR^���Α�*K�<���p������#���el���E�	��S�Y�o��e*�Cҙ����n$c�K_�t��S��0�I�S�R������'=���M��%���2R%�z]D�R�5�&��p��ጩ��/�H�0ә�p0"ig�d<Z�\=����Ox�����+����JS��3�Z�,:�������N��|�)�g�h�gd*T�"}(&xl�ik�>���/�}�
�H�e<��U��!����_���E��;����|�c����I�����I��p��篛�"Z�V9��-����Q�v����^
,w�g����曑�����G^�b��B
M�g�e~�%?����>st
:���uCySW���3�A	�W0������V~��/���x<��.��0<p!�p����߽��/�4d9�%�smt�Or��&����!��Կ�t��8ц./M^���?�+_��>pkC�HZ�ƣ
ov�M󩫾��y{X\��A4�e�Մczz���pGM�Q7��L�)�����Îr���xi�mM]od���y�mYY��]Þ�P�{�nHCT0j5�E��g08�$���8 2((
�(Ah��z��w�[���kx�Xk�:U�nwݺ�MGϯ>�N��׳�g=c��b}m	FC�p�p�Z7�����)�ا�l�� |Ȍ�DǗ*��v:�g�*������/���U���t����:
y��#G>��'�o�E �x�3i����</@
��(ɷ|�S��o����6Ts6'��Ǝ��,�
��ot��z��ͱo�UU��]χ��0_��Kl�mP�
�cv�C����5$	:t������&9u]SU)%Z���Y����T-ܛ��LY����Z���C�;x��U>��ky����[�@ �/p���(p����X_:���"�}߇Y8p���-��ņXضN����]��Zv����2<�L�q�{��=^��������
��^�B$�Df]HQ���:���o�-�O�E�Tl�z$Yr^ذ�z���*Hm[3x��Ck�5�P�[yQpz}�w��=��;ގ����Ŗ�� ! �iqj�4�L���;�{=u���.8|�Zo��1���s�AĕB�go�3����=���c�P�%HA��eee%��;���m��hL/����C�hFe��N5(�0Y,	s�X^[&�4:���\q�����[�A<$i��	u]�c�!�L�Sz�{&��Ñ�=ݩ������7\t��6�9��J�j�ڨN�l|���x��	i�Q[s�4�H�'�Ɛ۰����]���sF�!��B� o��6:��
)9��w��{���r��G��"�YA�%�p���YʣH2MY�\�-�(.X_���/�I�3�$�q	�v���u�NP�#l`�T�L��2�/�$��'����29�6���)%�^/Z�5��`@Qdi�9�N�Iq�n6�b����;�����;Ϩ4HB\im`8�QJ���F=t�2*KF���Tkn���B�3�5ue1�^%�S�*F�ֺ��S�����4"���'���K�R��K)q�E���!	���bfv�;o���K��YB�$T�E�R�5ݙ�Tؿ�V��`�� �aAx���cr��o^�01��
͜{/����H���=�3HW1�X���$Is�;�]GO��2�[w|�(�\�*O�d�a�`�Omý�g�I�����R"E�a���q"�:z��)��-��$'Kr��^��hX�n� *�l�a�3G�
���F�pD�� ;hcf�Q�5"P�B	�P(�Z��}�	�)U�v�$	�ީeh���(�Cnz���SH4��)��Ɍ:m�SI-B�"UH����iKa\M��B����	���@&�r��@z���D��p}p�oz�*T���W�s�J
�A���y�i�����!��2
:͵ZV�.�mu�!�2���*�r���e	y�#�S��28�ެ�8A⃒Hp�G��)������@f!I��,�(8uj�"��I�!t�.ڥ�B!F*�S����o�0��;���x-4��S���Yff;d���|=��jکF�%u�G�k�FlIiHA*Ӱ�ޫx=���k���є�Q;kPRQ�ƅlhE��JRGm�f�uc�k5��;���0��Ͻ���^��kɠ�(�8	�w;��IrM5�󬬬��k��D)$%<�T��DI�v۴�[��ʇh�Qʟ�]���謽V"�s�%9EZ�����j:]��R� �$T����R����Z3X끐�i-�<�.+F�!XG��[�3��W���\�d0�I��jSS[<JQ��eК�w�����5i���%�2h��Q���hd��&+`zߜ:^��f½5���
�U�q��bT��΢�$��rHߌ:!��"���ѩa/ؑ@;�����;�	1U9h�-�4E'	����J`}�s��X!^q���&eX�F�snBXzk'Py�����3�JH�BIH���� EBY��/�b�ܐL9�5*Tk��6X'a�6�7n��!D5�ҟ��۹a�BjPU� ���ހ�X�T���G8t� Zk�WV(���X�,G�
A�
O�j�s��>	~Kuۚ$5%R)�z%R�t�j8Zz��`��Ip̗@oا=�@%�R$�'Gk��)T�q�F��p��M�2�/�а��d�*2��T�V�C$��2*Co(q8��]�`���4�l'H �v$P)��xfj01�FA9T�53sst�f��2��xg!B���>��/�wA�������EA�w�"ǔ�jd)�W;���h�U�T	+++$J��0&�Jt���d�!�1()�R�>O�Rs�Gx쾗R��$����g"-(}�iN���U�n�9v�8�� !./�f)����R�[m�,�,G�����հ�Y
B:���(���b��{�J:+R�f�n�"��R�C�L2�0�ƨ��!����Q�5RA�H)}(Jk:i��*�kFQ\8��8�m�g���}�=�F"puͨ��u&��Y�5Tޢ�/�(�"�*YI�P�;h����ҬC�Qk�B���SVC6VNs���r�DX;X��ln�)�-���������Z���D)pW�`��9���TƑ$eYc�%I��[�AJ0^b(��E�jJ��uT��K6�m�.]l>=�r�V�hu�:g�%#c�B3{���~]3r�AU���ް�m�`�w`1(TL���OiJ��lj�Y`7J��n�pX[�\���z��Sx'�ʚ���>RB�
�LS�C�֗qՐ4W83��*4�Ō*D:m��2\ZG����i	hZ���-���7ґ	{���aI�5�Hq�cjKUY�P�,T��ZCmI$��8e]a��}�8����G���ʐ� DB<����o	oyӛx�3�9Vi�LS���z.9r���c�f&hj�����$�0V�ǉ�<f!o<:-��}����~���*�23�e8���2�H�	TU�4Kp������e�	���u�1���$�V����ŋ��ú�ٹ9dޡ4�~�����VN�-CD��Ұ�o����;���bn��6*@��,�T5�hR���]0bP�܃��^��k�,G
GYI���ʩ���0���Z�\X��b�K�����@�).�w�+�x�'N��fq�>n��v:Eb��I�Ι���%�!��E�✣����8z�w�X��$�	B+JS#��?��_�
�N�zܑ#G�5�J!�X[v��r�7"��Moz��Ϥ�m������+�%\���}&l�,>y�泟-�@7���xn��?͡�d\�Ћ�{e����C��������8�����a~�e/�QE�x)΃�J�{#���'������&Tp����{5��/���c������Y_]��
����>~��^ȣ����CV$l,���������əlJJ2$� ;�R�Ko%X
Y��%�5���]����^���7kk=:3��,a,)��n���u���5<����+���:��q��M��f�>��+�J�IxU^z� o8}�7�}�x���嶣�(�LPJѯG8%)M��_�uG�����@�*�sy$P/%o��7���<����
��}:Jqdq?_��M`�[�IaCu��� �����@�偪�PS/q�$�����*W|�#y���H���o��_�U@&S$SYFe�+�5<�G��gK5KK�1� e�Oj��e�-��mA�W(uo���y��,o�p��Y����|���[���8Ҽð4a�Q��k��x���emr"��(�(J�:m��i�AU�ӎ��\LYcd	�r���s��R6z#:y����tZ9�o��W�=��ݸo�=o�+6N,q�E��%)w/����Vgp�V��u�&k���0���Ŀ�>drއ��2����?�1,>�k�ݗ��?zӟr�oA"�U�І���V���@w���kW?��y��K��M7⑼�-o�Y�x&xH�d&+���|���҇_����̭_da4��@��|g�ޙA�g�c'�],)rf/8�__�i�W>���� Ѵ�gÍA(�'���>������[���iF��F���,�*�1E{�)'��ѕ�� <8c�i��֜>u~t��\u���G�m�;��}����w�%Iަ��Z�o��<�g�����9~�u|�_�Y���i�ز�ɒ��b�{�,a)�|&�+��і��1�	�����Y��~�y��1?�_`T	Bx���۾�[y����^�>��oƝX���k�N��t��U��^/LPFF��@���Y�v��]��)�����`iu�e��ox<����r�7=���+�����8 �9FH*��d����@��������`߾EVN,!\�x���8��?��_������O3�	8K@�V�vnAX�
O�AfC'��tn<��X�V��5��25���Ż�f���x痾���y��;�^~��<őC�9v�����?_�3��4��+o�+����H�6�KleC��T��(p�0�C!��ˀ8�a��~,n_�I���$em�G�J9����/�t�G���_���o��/�ȓ��1��C��ol�N4++�p��8��IO�ay�b��0��?�;C&5�N���3�s�~Xp��S���s���,�'���v������f����%�:q��_�8��O�$G���x�5���ۏ␡.�0�����7_�~��Gr��:�� Yf��v�ێE�	J���҇ճ��"pRBnc��V=�fp@W�|p q¡����5|�X\܇��ܶ��]�dt�%����5��7�/�e�����	����	����vP�=N�HB�(ڻ�᎘��x�O��y��RX��'����٨�52�3Òΰ�]UuI�ԴLMf*2c(jC�ttG���g��T�Nmi�-[���J�)Iꚢ�tF���hcP�!ڣ�y/Y ���qHI̭wp��"��ǡr��!0��>8J���u��"�(�Z2$��mT�@�^����"�A�.Bv�i�"�H��4^��']�*�eB-j��t�g�j��x��t
*��}F��@��X^`�\v�/�2P�.2��`[]>���\u����}�.2c�J��Z���b�4��K��!I9���y���%��b���]�f�bTr@k���p�f.)XlwBv<aX��P�L��jfküu$k�,
�"����tW�����o��\��u�ޞ��1�&3�J����kh���!fc��G�'a�2(�'7�ʎ�ՈthH���ɫ�b4"IG%r4@�����p@g4�UW��B�5��H�%�AE��g�����J�t�y�8dj�����G}�umq�Q�C����:O�x)�����(������b��t��a���5��$��<-�s��r��ZR�I�%q��9R�b�-G�!_b�X������>���*Ǔ9�v�I̖�YGj�5�PKaڹ����b=bԔF��2�L�*�%N�����)^fX��9�ٹ`,R�4%KۤI��9J�H��H�2U�j!t�RJ�x��ܿAW9V�8�`U(,4f±ފt��Y[u�25���[�t뚮�����-v�C�m��P��ՈjD}��+Z:��
F2o�Ո�hD0B;Gj�s�Γ{G������d6���2ki��Nm��*Z��9A*��F q��$��C�<m���<΅L}&W3]D��9A�	�,��hB2u�]Ș��1ɺ��fxr 56�/�ɜ'1���(LMa-x�M���"����#�F��!=�2Jj��M�R�MV6/�ʐ���XxJE�*	>�5b0MB�@�R�q���	�%��HEF.itF��
�V!C5n�@+�
!5^�X�0*��D	���O鈔��Ɂ,x�!H�Q2#�\jTt��2��mm!G�� ���
S����P ��He����
�xj�G%-Hf��)��:I��&K5Y��w5B�R�x+�.�ǉU̥�$B�Ƶlv�L����q��( E����c�a�"���Z��A����Sk���u�5�Z
F�S�`�U"���bZ�����dg��p��~���Y��Y�d*��DH�<�,:^���HlJ��`�4���:�3$h�QN"c���4[q��
nb�{gGsNmEȽ:��"�Y兴h����������b�k|]�n�RxT,p'D��*��m#�f�H)�rg�u��1Έ�<�(9�v���ӑ�8=p�`���3�����=�IB�$�m�p��[9hj'1��
�l�yv�Пb��������&k��ŕ'&��C��qLņTx!���VyБS&ށ���M<f�܉��oK&~bG��"/n Π
�#�Ɣ$"�G�4���*��b�W$F�딬N�LJ�MU��8�z����-�0��BZ��!|������8d��E^�>�άu�-EV(�\ ��CME%NTx9Y����x+�۹���{�>DlLN��*))		B$X!��"��"�h������-����V���ϧ��r��k}Nښ��|����ŏ��O8�j֔���&���:ԅ�ʼ�M�$�l���B��j�l�7Gk*�W�c�GƔ�!d1$��^�R!��A`e,(���	:�g����S�p�R�{�s?8��'hD��3���x�!����(ÍW_��Ƽ��	�fm�c"Ι\e�aL������:\kX���lX��*��I�������`h�]���j<.���#$��F���{�`&9�	5��Ͷ�AB�]M\�"IeN�@{	>�PfW_�U��G�۾��R8�C-�y��U�c��*N*Ǫ����"�@n���^ T�S��k�#&���sU�$�b %}�B�P�R������V�DPz6N!��,ԯ�lr��4��s�Iz�?p6���r.�M����7���C�D)�~ls1I�g(�(VѬ˔�J0:�V�JE�%*�3����91Х�)D�$pv9��ZZ,oב�	Tu;:�3+x��1��uzՈk)Q$�{Z�ж?$�5ZX��9w��e�Xjja�������L#�e�F�C�HX��CX�-�i��R�s��Uu�Ȫ��Hú��g$��J{��G�U�R;	�S&�i��sI�*�M� aI�O'�bUu�1C��8���>p^#�ҞZG]p�#q)�IP�\���ˋf���h������y�VA�Ӭ�N��jN�8������bY+�g��yʱ"c9O�g)C-�d ��{��)dg?8��2�	��@�BZTE>ܓ���-������\�������mp ?E���(�`�A)%Jh��L8aѺ�S;��&�����Ť�ބ�&Q�+!�'���mu9�k�	X.rV� :�v��X�	w���7�� )`n��Ds*S�(RN�
��rN}%��Ts^�>�}Q��aY)��Ť����V����un���)����V��v��V�R�Y�t�F�0��)���TR�d4�]|�z����Î�x��A�)� I����(�#�bM�ML�Vs�,���4��1s`�g3�sd�3���x*w_�����U�vs��b(`䡴`kF"m�:,������t:��!̆��p�7��j�����L��hۆ�b���>�\⮛>���/��'�_�Z~��ë�_�'/~���ǰq˻Q�/��*�Q9�E��k�U0JCiBh�(�bM��ͷ�H6D���̏�i�p�B"�5d5tDN&J�rs9�z[�q7���z��˒��\0BܵZs�K�Qf|�N�s�/��XN�w�O(�ߕC�[��c�"G�dك���f���6hQ�l����)����C�Y-xb!��[6�Xq�������O���ܻ���}���3�y?��Ȼx����/xſ}׺>��t�I��G߂�ks���C�\�Wa㘑��)%I�@O�7GY���8!�'ӃpA� T!�X7 ,<��I�-n_[��>O9����
�t�$+E��?�\~����o}����_���HԵ����m���v�&���LqV�(�=�s�uۜ>}���ؿ8ñۮ��|�#�şz2_�fF�ɻ*����'>
���dID  l`IDAT/�P����cmMC�l��%��5�a��zӐH��Ե�W;�j�S��l~�w^������7�	��������~�\*�u�x'�z���o;o�ا��?xm���]���?�Q~���䕟�,/��'yΟ��o���E�:q��G�5��GS\���qMP�q���a�]},.B�@��NG�q͏�0�����#���u�k��YJU`�`XY����_hw[��x ��(�O��F�
⡝ 4@˿�����'���p3)���a-'���̰������~��ph.8ȗ�<Nm΄�@�Q�"^���**���x��5Z�aȾ�zk�/�͑y�w~�ø|�G�_�}�����y��^�� ,<�!�'>;<��#J+�l��3�:��S�eB�R��Z�HL,
l��T	�J�����#r)��' ��o!��Ǔ<���?�	�گe�Xz别��I�_�(x�W��P<�j������>����9�c�S�u|3UF-�hR�D����%PT#%��� ���P-���.�����{����W�D������x[�к�2^�w�U���\߯8a4s�G������}���,_9�H�p�����Q�9q�0�$���sr4��^�̿�����|~0�cKK��Q��zf�;�3A�p���ٶ&A��B�%29�y*)&N�G�3Շ�gXV��Ux��<�����J������\�e��������|����;1���x�sX�N�GT1!�wed��[��H���ャ���w!RAgn6d���j6�� b�զ3ۥ:u77b��!�/St�l��
�~�[]�[o��n�a��3�;�n���ns'���9G�P��v���ĝ̲~ӝ���_f�#���x'��'��k~����*�9��[���#��3kK�2�;	5,�Rr)i��s5?�8��'"Q�� �H��K��x�8����`�o����/���^�����s_��T��ݞ��b4t���7�93^RI���B&?�B��X,�|D�A9�rj�Z(�֬=���tӍ�؟z���+��!��_�ç�s��]�e_��q���^j�|Ϳ8���b��1R��n�=~��鸚��"�mQ�_8.^�����>����5_��_�~����'�p~�������[x�7�+~�_^�3.:ȷ>�OǷ��	��]��������~�c��'}#���g����5�m��F�h4���'��ę8Ij4څ�4��&!K�ZS�Al�-s���Z��:���D|�&�������tHZ�m󬗽��"�Q���Ez�7*FUE:���[)��z_ hkNԼ���k,��}|��B��������&_skݧu����|c ��9y�\8�@"��_-CY=+"��z^"+Q.x�O�CC����Yd9��<�*�0p��}��Y�	j�Rl�������7<�*r�C3�.i~<�x��yL0a�{��1T���y$�Z8ā~�����,0��g��������q����}�C�O��QU)�<4oq�n�p�s��1�ڧ[f��|.?�Y��H�$���rb�j�pH+KIu�/P�vY�W�� ��h�ú�<�;�8~����r?�d�_��j@C�A'���靕X4�J��F�4�L��ʇ��|HOx���q_�\ph?�������->�;E5ׅV��;��>�hDb-�֔�0􆁵���9��vlK�+$��j��� pBa����ʀ�/��re�d��b����N:�.%��.�r���x$V�s�TIb��0�j:�$cD"FH1D��Y�����kH(j��4���������������[m�YJ�H3�̊�.����:�W���˘��.e�jf|�V�iaϐ0԰�
z���-)u�/3i���wX[1\Y*e����˯@�V9�g��3u��qç?��j�'|���3)�͐Q
C<��r���	���ٮ@4p��aLM�ݘ����=lb��z*|<gk!iu��u�]���rVVC��p�E����[���G��h0����=7��8��LnK5�gp<��)��^���e�{ӌ�n/lj�pxY�e04

|H	0�K��OcL�W?����à��C�z��.+�%Yg?�2�Ƕdp��^�}��9)���d��LDx�.���D@�e��Q[���1��0�2�0P%	�G#�p�$7/�R���|���`�d�yhw9�>`��������9mǍ�A�]#ǆ�0�\;��wDx7Φ�s�w�ԡ4�4K���ISr��󂀤H�[��[�ġ�9�O�`�l��U�O��� k+0����Il�������2�,^
���l��;��Z��`k�#�D��O���%P~�0M��I� u�k��P	�+y�B��_�[������#���]!U��x��^�o���`N���~�S󋜺�2��!t����=�	|�K�o{�/qsG��&���ޚ�3�-� \g��:�Ӂ�8a�U�R����&��*kP���)y�MRd�C�Ceaym��Q�Ae�ZJ1�n�i�گCE?��w�M��N�p��RZ�,1���u}̚c��tl曊}p��kK�Bp��!��8�f@�F'��Ë|JK�]x_Jn�%W>�kqC�����R]y5C�a�a�d^R\y1k�d��Wp��WQ=�_���o`��q{�4�)8��8g���"�kcmo��tШs��|�$HW�L�4�gP��?��UR�]PXkY�X��Z�#�O�0_���A�փr�����3:
]�6J��9���D�Ŏ*����������؛�s���j|����c��Ra6���zC��p��s�{?�K~�����d>�οr�$eYa����z^��o��x;���w�m�~?������{ķ|��`�4�\]��	N9�~�QB�։#�҄r�^[����=K]���QK�,4����\e,vfh'��*$�s�B��(� � ���i����`�"ɱP���O(B�a���9�+=h'���*	����?���������ûx����>�>~�y�EP���/���[x�?�}��<�w^Yu����x�;��_��7�oy#��_�"��)����6�yn�`'.*<!�r3VWL����(�­5�.�7�X+KtP	l���U!�'alE����4Ǘ5�T�v�^�>|�' ����n�bc��f��ΐ���j.�?B6p�ӫ���O�ί��:`R��A�3������k`��/�����Um��J	iR�u0�ABht�Ќ$�$L>:�ԮO凔��i�ѕ-擄6��?��Z��$�}�WƓ;K� q�]��P�v�W8験&?OÔ�k��!�����˃�rx.ه]�C���Mz�b(r趂�|;p��,�"�����@;%��zPnIG�4�0h}E��%�Ԍ�f$4C�C{o���H<˃5|��1�p�i��ZI^,�����<��Y]�`8�C�!�<-�˸�$v�!�}n�x�l*�,��<1�N�sڭ��c���i�q���󆷾�����u� �}��л�NF_�R���7���D������"�$;o%WX��M�hFzpK���rF�b��6�gfB ���
�jl�U��*RàN�4$ޒ9A�d0��d���X�%7��������O_��4k�k�?w�������G�;������������'\��?�3�Nʪ�D�?}�~�_pß�����Z����1��?e��Y�Z�?{����ڐ%!�*dk�Z�Z�(!��ӣ��KZ�x-��+��"m�.�Y���ޱ�:eĐ��Q9����/�+�����%P��Dp�I'T��q���w,�Xn�p|v��C����5��}�b�kj�h��`�4ݼM}�8?�]��=����G>�W~�7���|���������|'W-f5hY�3��B�6��D��TexK�~pW0�N�Gkl�!C.Ӕ�x9 m�<##FԲi�ʑZеD��Cҗ󁓛�!O�C�X�T���������Q�Ƿ?��x����y~㻞������;�;�/��Q��������;��W~�7���ɴ��������������o�6�{�K���|������� ��:�<��Ā��@�
-�%چw\/4M#�B\��v�`˒}�3tg��jS,.0�`�
����k�E��̩�V�#
�a}=VH}%q~#���C�#�Ʀ%�L�U�Y��G<����so�>�QA���{�o��w0#���]ą��",��Q�|��o��_�J��������$��D�������&�JM�B��F�F&A
85��/ ��b�H�q���:ݰV=ك�Rj��
��>�'���� :B�T R#B���V����l�����r��k}\M�,Cq��Ŝ�\"5s+��*�w��V�Z8X�\P����ZY��*f��������1�4��4b"41Z��qTJz$V(�Wט�?�zY�����_\;�7��o�N�pç>�h}�\C^� 	�4=�7p�`Gmꃞ�R�+�ZJF�aF��k'����_�Ex�5��e�ið��+������/y	�|�A��d<�G��L W�r�a7�B�tWO��-s8��ġ������@�BU����50SY�j�P�L�����y��2E�c�#LY���X��O�p�>F�M�rj��"��������"&M�b26|�M ���X�aEg0�KI���Q��V!�A!`���.sJs�hsHe<da!h٫�+�Ԃ�4tjϜ��S���q� #ä�$1*�^%�J\H �8�ǘF�H(e��)�3�m�!�[9�-�2������'t�q#�Goc���?�Q���J�3q<�8�5�7��&p�3��Q�h��s����w���.��-,¨d��/?�Ы���W\��sA��<�	��cme���VUqQ����p��R���TD��*c�#DH�D�Є���Y���*��O�>��07�����k���(��88#8� �%\��cԮ��9F���/D�Hj����Ѣ���ȏ��2� ��[]a^*�$-Z8��sɾ9l�C��U3��>N��B1pY�G�a�BeX�9�0��TBG�$B`��j<�� EaqV�CyB��H�(XK4�yA�� ��n�%����G>��}ɯ�`�ဿy���囸da�L���U0���l���y%;�x�Ʃ�8b�b�y�%��dޑyG��G�yڮ�5p�N��[�
7~�N�_�u^�����Iƅ��-��˟�<dm��C6�#��	���%��_[r$Í>Ԗzf?�R���!�����.& k<�Z�7!��cI
e5 /:�|�3G��B���3y�O��I��䱗��<�;hK���{t�I�l�K(B��$�czxl�K�1Z��`C�q���{�5�&Tplp�X�=8�v��Y����)�Q=@
GW��>*��u����h�>����~d�Loȱ׾���ǟ��X���8�~��<��h��;R���B��c�ƽf����>$_��!4!ߔ��ʒ$/-Cc8���-�!r	�6C>T����9?���7x��^�|�#��c?�	>���઼Ky|��,�:acP�8)Bj��`�ɘP�z�yٛ1��v|J�|�g�f_E���K�f�f���7�/���~�����ؿ�ƕyN{4d!ST로ai!�����]�ZPII�&�@B&��WM.����( �����a9D&�$� R���}�O��o���x�K���y�/�+���q��������s�-+Q��BF2ЅT��y�-���#7k���(h��x\5"�9~����_z!����'�bA+
ﹸۡ��N>�o�����|5�cJ�b�@��	�=b2�#�6c}�7�z��3�.�,/!fy�/����������W}�������Y">�����+~�y<�+.p�Y/�.�I2�ڝ�<P�xR�_$b���P���	�ƵB�R��+�|�N���t�W9��H���F�`VIB�Ň<�I��%�D��Jz�c�����EJz�"J�:��>�i���0 ���<�vm>�yǻo�3_�M/�.�\�g��_*y���χ�|�l�E�$%����!���c���4�+�QyB���a	��#G)�
A�a0곘�\���G�"]9�W�g.���%Z��S�ɖNrU;�0}�/�"�>'ш�	���s)'Bڜ8��eSj!���4��]��X^�QYD�eWm��7����}����'��u�;~�+��������[$&jՃ�Q��,�5�8)��
0j$k1���y�#Rq��\��OrD�|��V�+�m��n8~�p��<��+�[[H�-dX�������1�;�6}pc˵£�ɚ���}`����$o����Go��?�ͼ�7��$�|�?p��O1P����Q�&Q>p���q^����u�3�yB:S+mp��T�H�Ɠ�5��HZв��C�2�����2�XȆ#����]c�Do]��M�EH���v��;�>�� 4����˿ʫ���??�,�����k�'x��q��G���ٟ�]�����G��T<�K�󖖫���A:K�'���Dv_i�8�G�@�AW+I�B$�Hi�IF/I�'�U["�E��|T�l�+��,�zfVj�/��/���y�Ͽ�=�$����f�v�M(3�8��਩�g���#��bSL��w!ǯ���LeqƓ�m��]D������ɒ����-�w�w|x�����Du.�7�BɠY��\�/���'��袢.8�'�Б[EWJRkq�ud5$Gb����P{���zM��ܧx��H����E�&�)��1���ϕ
�O���l�T$ќ>}�,�u�C���Ǿ���|��ב�s��
��O��\1��$�v��P2b�*,��P��%y��}��Vn�ID�A��I��ʑ���L�:K�=�	2��Gp�L��mo㖿~;�g>�ʧ>��y�lmh׎���*�A���jc�MN�Ŧ���F�Y�*�*=΁��5���T�X�wX�s��ǷJk�,�{:�0Uh��C�)G�؅�^�},&��-�Q��H��#r4Ta���"Ih��V-4����~�Q]RaHQ̴: b�^٬��D�Q?{E����^�h̙���Pd���9�TH7��5iƑ����%��y�Gm.O檊d8 �u�	�1Qj�GZ(���3r����7vP����B{Ca��0S[��%���)G����!��Q�^��$��Ъ�t�>u��
�zHjj2��|�SM�N��$~>���@m(�"�0`|X{��h���B�3T{��;K63Ckv��}ig2���I�=��q�KI1�|Д�ba�TJlP�%|Y�� �E�-#[ѳ#�͐A=�b�����:SF����	���Z��IEE��BcH|p$�3\0�e֑X�V��DF������f�@3�m
;"魐�/1Ð�[-.[��¢E�Ԥ�!/��-�������.��uk��+��^Bb�#'�#|�{1u	Q����u4�v@<B�� EH��.ZA��A(Io�gX�K�1��}�i*����
�&�'����~B��1//"L!am�d��|�f�ȸM� p+W6½��fj��W��L��ێe%�J�YP֒��2���&ߑD
A"�>�B��p҂�(ob�{���o}�"D�H�H7�Ҽ��3��V��D��D�B��3x_�0xze��(j��^�� Z߅s%�H��OO�X�5��ה>�9ý�l�ӥG"M���_��F�a���y?�_Y�����LYc�*h��Sy�x��-����#mB��K7��}�&�֘��Ŏ�q�I���T��Jj�q(����&�H�0����+/1�HR���2!U)Z�R�`$F+ȳ.*�#-�^� ������U����J"5���{�PDV'8�P+<q���2A��k��E	���e��X�C�PZ�tJ��B���E�
:�Y�v�D%���Jd%�|J.S
�,q8�v�:��%�cK��-���T��,:�!�N�.�"��P	2k:���1�'x;�J�ro�م�,�hSs����dy���c��+���ur,:��<ū�|�5�e�J��nHm�(JW�Ң$8�18&фp���(	���CnA��hQE/1��5gfT�(e�Uņ�fr��T�4Yڡ�u.��R���`+<��3�P
O{f�!CZ�����L�0W��3�����2A
����bZ��xo��(eIO�y�P$�V"��y��;���[�V���5�%y[!�,��A�8p��z�U��#��!�`��Zo�"��j��7~�ݧ��y<c�X��FJJ<�de�ǅqqږ4^��dR�,t.84��m`�`h*��Ћ�oCc�ꊪ��F��~�dy��.2V6z,,
��I0�WUE�4�\����k�uE�$���$ɰ�3���op�`���`�v����1[�fLEe����Rې��Z���k��j���:�L��yNU�6�i$KR����!N@�����gv~�C��e����Qtg(Z-����%VK��+�!��jҋ--D
;��M����>���QI����W5#)�s�x����p4dPQJs��)(�x2S�~�(�Hѭ��р�3�A:J7�6#LUR�5��)MMmC�LMY׌̙��kJSR���R������,u�I��r�<%�v(��G�iJ�(H�ɭu�7�S'�B��� ;FJ��y�79���U���r�p8D�F�I�X�c�&��#�f�+���B��T� 2A�%n�g�7���c#�gmR�,v��JI7�e~f���ţX_D�`,UK�r�?�\|5"ϳ FyK��>�3�52KhͶ@IP���\�4�I)�B����;7o�/�X*Y;6����kF%�&�p�ЅX�C9=^�n����i�{�������jֆ%Ck��`X;j/1>$���T�K"xC�X%�l͸ ��$"�٨\0����+ش`�%�Q: A��F)A�j�$�[A��6��S�Q�������V=6�z� �(d�P�Bf
�|N2�"I��|��[]�K�M�"�Ԡ�J
�,ecTAe��I��aI�$�r\=
��8�bGm�,�Y�Ȉ��"�o)&��	!�tf�.̣������fUJN{�i�Yr�d-'kϠ��ٸnk+N�گ)Ɋ�;�kR�T;��p�m���Ʋ�`�ŗ@�ͱ�A�Ђ4O0��#׾�\�L*��G�eR=�HHV��b��M��I��$&6[�Ė'��T�1���6k���\�L.���:�sϥ�99��-_p�v>���(#)�T�@w��.`�ZFyJz`b��i3b��%�=�ӂ��Њ�RlhA_+z����zZ��_8�Ĩ�e#-X�}]p��5t�J��˶���xg|�_��y:�ƕu��~q�~�a��J�E�Io9�B[��S6�K.�U)��V�����%KHNXϨ��nk��2\p��Н���^�7�Ǹ�4�a�j7ק����N���_�Ao��@�AJ����[���O��-�п�ap�V���@������կ��[������F_L��5F��x�UKٸu5Љ��Yd��.���^Q�%�\��7}��W\čk��C���o'�?��t��_��Ҕ�F�UW�>���}~������JRZ�:M��3��qM�����6/���l���7�Σ��<II�mn��fN���oz�W�=�|����<����{����Ri\U���t�ND������m���y��iFQ���c!���P���^`�fiT�gmfE�uP�97��"/��_xͫ��˸�1����*ƃ�4ê������W��oz����ՓK��#1�\j�^cI��l��i�:"j�*[��&?�>�� �����ɾyn:y���������~Ǔ����I^�淒���CP
����~�\v�e�w�(�</��a�Lv�=�Aa��hL�]ȍ�ފ�7�ٟ�?�c���$��FX.��7��r�_�=b�����Ut��1��$�������68��<�N#O��u_�P�|����>.��Jn]:EՐN�Mo�� �5��u<�9�����p���� �5y^����q��!h�8� :����<̷SVNo`�'I��<��i�󟸎'�W#�#M���)Z���/�*���?���?|����;o��vQ�Քu�I�s!SJ�3~qt�X�t{�Ep�߾]z0
j�07;ω[���1�Қ�~8��9���>���������]|Lv�����9�o?���?����[n���{�++$��f���k�dyߍ�]D_�R���%���ʰ^�pݜ�y}���E��?{#�����ң5;���*$	�Y���*�w�?��#�_��R�A������o���:�|Y�ɐL���y��^ƕ�&<�a�$�	�����K�f�����!p��_ �Y��N��o�Kd������Sd��YZPds|�������QO\vS���m;�L$*���->������/b�KS��������~�'ǚT-�IRUPU�,m���!^�[�� ��6yc���$Q�����7)�=�k/0�TÆ��S0��m����s�CoX"-�:�.��C��K/�9���gA����p����C'���8�2ݻ7�0���pe�W^��/�m��mo�K7�N�� 5��Py�bVp��I��}ܑC����K)��!$\qa P�7���x�3~ �FX8j!(�9����n���Zk�$�Z�[+7��:$i���ۀ����0�j@�����jK9
�,!�����:	��!:S�vfY]�蔪�����u�x�`��� o��H7���,����3�s�z�A��E�)�`�`7֐*����q����<E"ی��!X<0�s~�G��'<!h�������� @'�i=&����N;�$ D�q�k:2�P���|�S��U��;� E��F%���&��!^*\��ϵ��Vװ�e����c+�Jq�!rA���,�h�UW\ĩ;�2P�p��Y�(�(o�r�giKM�? ��=q���9r�w�$�T�Fh���Y��<�s��|�_�O�~��4���{;�Rm�?wgl���">�{��!��u'���P�����H{�.��t�k/|����o�/����-�Ύ�B'�����ucpL0$X�
Ap;_��VL����o�\:^���	�J�-�
M~Kr13)8x;�@��17/���7[`���p�҇{���D�F�-�b�w��$ee�Rs��;������4Mq��n�{���A�����"ƅ�Bt��CUU�o9��ƈ[$³5/�l��B�����-l`r�M|ܲM�P�^��#�k���������a=+z	B����i��/$�#؝�85����'�qc�ٺmr��[<wă�X�ڠƉ��BE�C=��\�O�,b�&h|7�c�yʡ�g�iRR�|�U�x�sB��ނ"�j�I��.Ps�����_�1gW�L`s�M@�0B�g-x��XR%Te/��`����MM3go��f�&�����ԅ8��F6&��@b#� Y#���Bܐ_>���l-��Op��K�E^�x�pB��	��
'U<j��YʐW�X�*�rȪ�C?�Ӵ�lB����[%P
(�b�����epP	Aq����h������mN�**�$9���!��'{j�qRc�d$$�����-�iˊp/ab�$B;&䐅A)5~h22�u�5��,ؑ@���1���'I�T	 ��͜?�mD�f�d���>���C�KO���H���"�N6B�����|���c>�p�{l"�������~t�w"$�nJ9z&�*$s����4!�LlJ'"BD���5����ij�}�,Rx-�C�e��F�m�{�t�W�/�M�0��E�����Y��@`�R�����M�qq�s�\�"79h�E'����*����Cz�F"l�ѳ�O(V������A��4"�w��嬨nϭᐡ�@(0�~���m��<̓aǍ@���5M����x�͊��/�S�w{�Iigi��l��LXO��0�%7_��?��Mom����W�=6|(� R�lȐ ����GG2���<V	j!BFH�ƞN�RHj!�c�?#��t!4�`^q�1���;�r�ɝ 	)����f@H�.��R�D��Dzb����3v$�A[|-�q�z,PW�8���g߉������cO3q�c*E�⿇��o��Υm3��L�Ṉf���Sx�A8�T'+�ś͠��٩o��k��HT;��5yx�@�ɇ��g�@��E�c�q�<��󖯚��s��)S߬�LP�L(Ӷ<N��b��&�*̡�1gk8�潋hҋ��^��!zb��p!0��C����X���5Yk7�ѬOA��R�=cb$l�kH�>�P��}����2p�(��E��Xք5(q�6�C��ԏ���ϭ�|}�{��&�Ć�MX『%։��ZHL|�҅��1�&4*F�g�2d�ʆ�zPѸzf/�
�)8.�kd,��}PT�_�@c��w1���j�:�V��A��6�-���[C����y��kP.��O:ݚ�P3�"$��[�K�D�s��Y���1Uf���ѭ�Q�!V%dZ$���8Q�����+C%9ޅG���@��y���g#иN�����*Q!B�K/�db�$��ĳ��=���/�zv��&O��ق�u��oy<͵4]ვ3��v�r��C�,�r����O�c��f��)N(���l���;<��m��4;���I�[v,���\�e�7>g3��v ��a"c��ɱ��5����}�!�m�j�>07�M4
."�L�X�gbSq����`�{Cimu�b�4�
GmJn��f���<��������A�Wh��	B��YM������ߝKk&��GV�m�����KlL��7��7�XFk�M������#DPia�� ����xj�F���Z�u6hҭkp��v��C�5&$ng���`��m0&҉�JC��6��&��}&��Ha��QAd��!��ȇ�4�o���"��|�4��e���w~���k,
a���z��Dw1�S��rT�� �4�5�/���/J)���-�k�4m��޵��8���+����/@)���! ����<�)8cY:y
g,y���t� �!W_�&&����1�ǜ|�c�\�4��ژ�ډ���N@�~��v��~%�*��SOS*ԫ͵Z���7n��&���9nh[��B�"*�����D;�7����t��&)��}�>��l��9 x�l�۷Mn?�~S{�y��M�	��$/
jkHҔ'~㓘��E��N�i���
A
@��O���Y��x�9u�ԣ�45ͼz�e��4M=�[�������ޗe�_��������Y�y�k�=��<�67���b��Mmkۿ-#�V�[[�Z��gs������6�$\Ih�>�w����5�����_�׺�~ۿ���.����K/��?~�7���1�4M�x�eY���vo;���vt�[ZZ��C�}Tk���6���(���K��[�����ѣ�Z-���~���o�u�{G�%MS�<� ���޷bR �6���M|���v6�Q��V�]�o��"��K6��O��'�����\�Վ��E��ܶ��b���܆��O�����@#��_���Q�5���\}�ռ�կ汏}����~��|��}BfffX[[#��&�$x�G���r�p6}��Ç?j������ԩSE�p8��/dyy�p�ײ��� L�y�c�{�D���x��T0A\q��;��c�~�x^m��!0&�\��Dx��]pV��A����_i�<cJB��w���>��?~|L Y�Q�%B��۷z��������Hk]��N�Bk����]vǎc0p�m����?��������-:��%�����k�3�xM�}���n��r����'�q;���u4���c�W�g�~�=���}��ol?��p�wPUJ)�ּ��/�'~�'8q��V=�e!4��jW7�#���}�#y�w�y@���<Ǐ`ff�����\s�5<���ۿ�۹��+��>رӽob;�a��'cN����]�?�F\�	��F1t;�Z���!BB�3�1�r��9(QD���	x�	����l��M������H�y|��7\���>�����zcEP�ۥ���k�֤i�`0�ȑ#���ۏy�Ӫ��}��|χ��^k�R�����RJ?33��4����>�,y�E1ާ��`nە:g�I�IT�z�[[2�,�P������%c��Z:фG��o�ִ滨`��ߋ����{�����׻�v����j���}������m���n�Ϸ�5� ~~~�~qqѧi��<�I�x�+�<�1??���g?���t�S�q�K�d�iO{�������Ǐ��tHӔ�hDUU,//�gE��Y�����Q-IR�h��U��H�H�^���2�e����;B-x���!�B)���/��!pBv!-"X�æ	�>q�HLb2zvA��!M���6~�уH � M�5�6�3)�߲�ᾚ{���ͳiR�h��b_���voؾ�}���>BVWWB���L]הeH�9;;K��E��W_}�W^yݶ���۴���+���[�٤(�� ���v���Zk�Z������W*�Y����K���	=ìИ�D�j���y%s�t�J���&�!�PxH|�e>ɤOR�u�|�e>+r�e�O�ԧ��*	n�BGwU��:�J�a������g�T�H��U"}���NZ^�,p�� ^����k��Zw�V�Ro�nB�1i��������Z+��E��<�B�$�WJ�~����Nogkgl�l��G������74'\\\�����m���MJ��<�� �֩O�܃�Rj�$��z����^	E�@|��C�[ٌO��W"��Z�|��|"�3^�xb���kI<N�vs��i��֓�	ğ�p�YҊ�7Ǔ^�$�i�{-�(Ƈ�"\g���i��J7�C�򒎇v�?����$�I��N�3�&��?����B���UeY^�����vTM��n{�����������ؖc�ٕ��2��H�]�n���> �VNmJ�	�$�zk�X�R"E�߁CG�Z�B��CKO�B�^�@���Ţ��28f[8�E�B�\K%ޖ8�c�)ʷ�_�7_!���@6�
�_�?V8�78�{����a��	���E^$(��Ϣf?/Z�V�����v{,�	!Ȳ�D��q��a�?���������~������g��{Vl��Zr��ѯ���֢(D�)���o��]�E�|�	���;ڧy�ZRm6�	S)���E��4>!�J&�����L}&�OD�>��S�����D�k�O���P>�ʧ�>!�9]_�Y���gJ�L�S՜GxM������k��g2�k5�O(�|������r��^G=o&7�'�'�&�)Y�n��T���iD�N��ݮWJy�Ԙ��SoB�$I���<��}�{�3w�9�v���sn���_������io{�۞�����Z�X�0��oGo��;m;[�����<����������vvv`m�t����?���y�䁃VVz�P��A�x6:I�I��� ��+�@��j�$�T�0B�\¦����LB�\�/�q�Q"R�h�Tu�mP�E	E�t���4)�6�O[��\I]W�D����zGP��!�7נb��|���lll���W^y��M�$�}�݋J�Y�s�{��n�}L�����b�1�|nZ,��֦�j���'~�'�'���.�b�ӹc|�s��	��9�����ͳ���'>�_����|�Ӭ���$	��,�������d
���w��"�t;,.b������E��y;J�e����s����O�=K�(>�ῧ��XW��9�Y\8@�=�֚���b�����q�$�;��dn�0E>CU���WX^����% fg��0w��<B��uV֎��rcL������.��t�z�>}�SK���H���<��,�\��ڲ��cii��S��JA����O�^n��n^���?��O}�S��F�2�.1%�]�.<��/_w���"��qǍ�zH����Z3��\���qu�[o�(ibɋy:���~Py`�v�]w�"TUˋ.��*����7����q�V�@*f���;�8�h���ll��;C�=������<�f����QN/������\I'�Yɨw�N��h4bvf?��9IHbV���r���%��t:t�d������{k�z�����hu��\Z<��O-������{m}L\ѳ>���",�.��+Nqw-^��{���H��V�)n�8]�;�;,�[�~�����&'�9��93s���&�&�	����^7��N�ŝ�S(�x{��C]���/�/uO�I(����*�e<��0����g�$��d�m��mόM5��>P �I�
A�N��-I͉ʿ��k4��ζS�n}ɽ؅��'�>�K_F\6+Ctx�-%�)a�[F�s�@�����6ԣi��S^����V�D�3�z����C�m�}�P�MQ�6��s㡜s��Ѱм�α�KQl�{	�30p۱�){]Q����������ju���d!�B��U�nUL�K��F�e��i�U��uA��׭؍蝄A�o{� W,u�Ū2�3$u}�)�_U�{8�9a��!���㔈3������Y��9��w�Tk�W��h��o
�m��t�@6Uu��%��f-l'��;p�O,�a�8�=��R,#���Hb�_'kj��)���;�l7i�~�J�lp��M�P�zu2X� �����Â�$[����y(yf'���߻�����1�}pP�t�b��u_�es#�"wR�dX���q[�s�BF�˃V\ć3_w+�0�x��H��@���w)�+�܋�B�h1��L���=M		� ���{��(*|n[��[-}�����Ӫ/�y��귏5$���a������h(>L5�+���*j�Y��<J�U��x.�x�EvNϒe8��1'!j -�/���[X/y���hR�H�s��mΉQ���Є�/eYM+0�9BO�@%�v%�7�G����&�$"�h77?��Jn���nl���h��d��e:�zd}wy�
�Y�f�W�S86gR �a��#��������3�)yQ�ŗ:nH�(g#h�q�!���G2Ԟ!����X�{�<s}�D�LZx��{?e_��)��z1���2�!i+�G�qon����M���@��C����O�⎄FM0�Tn�ѴX��g�C]�����~�q�|�d�V%ʣ����ᨉO����Pr��H��I�	S**��T5�_i~|�5h ��tV���u64�`n���kiezp����>��TA|�7��\��<��&�uҘ�žO��\0�:~�^�A�G�ޖl%-�E�"@�?�h���
Φ�a��to�n8����WG��0tߍ܍��6�� Y��d�~��,מ���=���m����v'Q� �O��u�?���1w�����
�U��G��.��׃���;��]��vؙ�F����x:O]�[���'�V+!<�	A4U�J���h�-VL,��]m]Ȇ�,�0�ƧN�������!�'��y2짽}ǆ�O�.��c�H�UE^�Ǟ�u �D"\"�9�Hm΢�3�U
���Y�%�	�	u�'�ш�ū�g���W�JH�k���T~�M�/�J3��ĀR%��|�c/|,��ڻ^z��`���M|�(<�Ԫ����~�U'dx��í%�����w3.6�b�R:Z��nr��HÖ�+,/K(�x�E����&AN��&�+�l3-�G������ᕗ�ȉ�;��..[�R!���l����[_����tL__��Q�$���q�H�[x@wk��uT�^�0���P<�H+N_������e߂�Ba�d��LH��$���ng�8�ƹw����d���ń��Ϳs	�H=� ~��l�(T�g(}���oY_|�/���.�G3H1Uʷ7E����P���s��\>�l(��qXk?#�VjW=H��Xsd��q�o�8�/1���눫�~��'�������zW��Aʜ�!D��/����lP��U0�ީ�^߮�c��絅^�g_�my�����wVh�s��w�&��?JI�����/����v���/mhzT�o7�a^b���{��/�V�#�������v��oǜ(yWÍ���A�2�6�8�aϊ8����q�5b�{q,��~l�X�l�2'��������&Y�1�gֆ=�K���G֮o��ʠ4]3
Q陏�J!�[�SF�(�,4��yw��}�1���"W�k%۴w��� ����b��� _f����VMw�x���A�t��=|e��	�_>�e�J�lJv�b����p�o�Q��Q�}�3pX-F�c����8�E
���a�e��i4�}�{�z� ���FH(�9�`��s.��2�xqV��t�k��\���������i�C��-c��:��g?r��L�?4�z���~��U��P�{bE������~ށլ^}��a��;�o	!:�6�a����O`X�s5���y�O���^��Ҥ�{%��7�k(lc$������w��?��_^�坡�@5���2^���<�M০
x�f��o�ɱ+��d�r�����S5X��;��;�~�T���Ѿ�����6���Hߔ�b|DgrM���"��B
��cg��s�`A¦l��3�`.��.�Usq
~�&�{)����C{��O M9DH��竐O�ȷJFQ���$������S"��Ţ��7&��_�8�ĔX��ހ1�A��?�S�JJ#q�Ȫ��>K_H���LH�Rj��J�%��I������c]V��)^3ȩ�κҙ��=��9�!.�p�Єz���x9v��|ĉy*U-�mX�U��T.6�1ǀ����77��ϗW�Y@("?cO���z�@����n�h��<�:M:ΪzS�6so!����"M� i|%y�G͉�f�U�;f^�nhO<�d��?@������x@��\����&�A�R�d̖	<h�1/�@��?�e���]�8}�� `h� K
ESL8�HJH&�"�_|J1���ǟ��_.���`J�N��%��{�yټ#/q�N}��/���fi�]��rX��E(� �%�o��*���Jp�^�b��VT�� ,%�)*5
�AL A���e� [�%�T`�.)F~=L�baU���{��W�T�_b��Dx��WJ>J[����:��)D8�JP"���ܓE!�K'xm���kt���Z����Y��<V^���H�%^���@��'b���V���i� ��o�ޫm�T�I�a :$�VP��ǵe��R�XP�W-z�-��(�H�>����p�8K����0�b�zS�,��Y/�t	����l�g*a��_��%[-Ak)��.���g���J[P���m�]1��V�<��$M���ij}M�T)P�/1W3\�%el��y?L.5���"N�"QHF
���������k&��īn4T��4C�%��U�C�#���QXl�܂$�*�P $��K��z�a=x��f8�`��v�Xc,b�L_�Y��Me�Av=�@.ð`}띵;����n���!|�R���|Mb;o�b�^���|]��9�e�+�C|+(Q6V������
qʏR�i�L=�Ũe�z ���q!�D�+�
f#�[���9��XV��~���/��]�}��E
��r�h� 4�Z��&꨻���Y�ϨH9D�0��Nn��<L�M;�-7M��s�.;Ѫ4)(��?���
"3��m��	��%Vԉ���z�:`n]{Esx$��-i�/�ֈ��JWK`f�O��>{rC,mMD/XD��L�Ҩ��K���M�E]Q�/��+�K
0j���Snq���F�ZQ�\	l��
�F��/7>p	��Ge�g=� �+��I6�(�\~��*�7�Pǵ+!ej���jP�!-��yf����1^���q�{LNj_CTn�1��0���.߸~�	�~U.��n���L��1���K�(��W1�4���軕�����v�F�n��-�;������a�٥�3���=�A���{����x�vs��qu'�\3�O �V^ؖ��R�����6�$��5�2�-ubj>��;rmr�]�_t1j�B�z���*.�H�j���?�4?
��B'����>�s�����!!ԯ�ð2�u�?k���^R�Fd1�U�&�~���{����.��_ ��%�-�l%�ڟ����8�6.AB�`9>��,�����"��SA�_��X�Ct��p���y�(��� �����:a�2NH(H(��=ir"7�D�RC�<-��k��p���]�x�:ẍ́�\p���}�^�Q`O�\��*�k�F�ȫ��ѹE>�W����7��r����$�0}@��5���Q�q�]iސN8�T�2$� Ga�)��,�L�?I 2YW��k:�tGX0b��$���0��U?i���uI����ts��yq'y���c����7N�G�18#XF.��o��*1j"�%�Ҁ����jC��J!a�4��� 	�g�Z�P?�}��m��^�J�� �'��wzYġ2X��e�_���۸���r¼�$)���$h3�/*Ła��ab�a1:��r�R�^Ѯke�@��H�u��jȶ��N>0i��h�U�esh���ek�t��g���mw�o>�(�W��rż�z�Q�Tr��������T�S̕!CP�n�!s�0w|P{�*�P���4Ǚ/�f���[��<��f�Q��wS��R�d�W:*z���%~e��/���-�Wqn��.8�bu�u,�wo��cVam�|ˎ-uB$���Oh/M��l�a�;�;���^VC)�^��`�]������Q�����|�U�Hw{�[�j��~����dD'�Mg���pM7�ZV؆ƺI=+�E�$���H?����K�}'���d����x����&m��b$���B�9߇�qSm
��@:وz��O/�$�맺��2�����O�>��;��Y���³�_�"�v��|k�{  ��KW��2�K�j��O��P<�a���ͧ���������?�+�I S�"�f;���ɂ^&������&\�6;m4J胲b��Ic*yM��R!&��rO��q�z���J ���-�����H|JF�����c��k�����"�a:�a�u�=�F�$�Q�$:1�ϸ�zjv�:(�ƕ�"&�}?L��r��SG!)R�H����P57�d��I�'Ֆh/��@�P�]����S���]���hr>����N5�=]ѥV�?�Qϴ=�w>�Ѿ�jW��Zӂ
��b�׈�� |������xǍ��Ri�@�¶�d�O���#�S���Y�^�E�FР�%mf�/�SSK�hV�]z��Ȓ̮G�෾f���q����e,ee6�*�ۺb��w+�e�İW�,�}�z���V�f4��Wh�+M� ��m�����ʺZ�9�,l��E�����X�H{x(�`Y{�Fn*۲KbF5��C����is�es�9]��&	����`W��;7�N���߽��J��M�1,��|�@#g��(�c�%�Q�4!��u�W��Gؖ������9exn��u��z$�����g�w���&���ĵ0$��y�V{���B8٩-�c�0c�q���u�ǆbF�����G��p�nԆ�R�|kZ�"%T�ə��Jp�čAZcK�NQ˥��4{����y�܊^�S����z}�᳦1�?�b����"�j$c�b��o2��O(��r��I�I�y,�!�X#B�:���}NW��6q~'"�.(.�/��A�Iw{h��i"1���;�>�&=�N�C���g68b�������j���ģ���;�@%����鍵䕚���r������ ��"^�Ϥv�����l*���� ��Ͽ�ǵ����;��g�N����̷�'<�ob(��@�K\�G?q�Ƿ�������}��:4�-�IU�8�,��v��_����g.-ca9�=0%J�$�g�U+�,�ࡀ)�}�EJ�oy�bz7�)*|l��~A�B#A6Xo�����4�PXYkL�XGH'���T�Jh�:f�0�M5PdJ<:���=8w�)&TI�S,���X�R.F���c��>,�#Vj�|'lq���3˫4ͦ:�x�����GH+Z�؎�K��1D��`*��n��C�^�id+�ߌ3�/Q�5F��.�eea��|ca������0��'��K];5y��6;�QKk�K�	�]0�+[Y.	`�A�Qɪ@�+i��4�#��"r���\Rǵe�n<4�ox�$byy9+Q�9�i��>��g,-�C�Ņ���@���&�o�����?��d���4|Jp]ř�����cB!�~��u���y���%	E�����f�֑f��=����\�(S#Bǵ*��4K:����9*~�DĴz-���:I�����W��գ�>��a�q\�#�\h��1�� �~13̴|)�&��u�YV�+�S��b���󟗕�jZK$ُ$Q@���"���g_Zt\��<=�Pk���S2�8�5����Y����5(��)���O�
��QX����x �L�~�fn<�Q8���T��lR(���K��������� X��{ ��.�������7����<��>�ϛQ�ou1� ��AJh��5������cl����"��u��U����www�����7�)���b���0��'�w��;Wˇ����D�"��bч҈���R���>"ZS�(�~�z~C��ɉ�7�+=���� :�`��~0U²=��7�39AA\��c?�P��	#Ax�Cq�����w6K�_�&�H��wD' ���=�'�I}<�?��P�#
�a�K��	�N�
x<ω�Zp�dkkkC����Oc���c˹�)�����u�V	��t!^�� ����Z���͍nL�{����@��kO��ك��;�������8�e}�oC<����:FL�% ��FFI)y��o�jW��~u����Wθ���6�,�|Ҷ@_ǡ��g�%�e�һFf�D�����M��9�Hp��d%'㕕���"���K�Դ�����[/6�w+�ܧ��s���k�+����;M�x�6��.�.l�ֳ��;$t��;99	u����T?�շ�{��'H�3�&It���Z�<^K�c����Fߠp��=7z�ФW��{�+=�3
��M��"�.J�o�Ც#��
!�#x	���x��X�����4��2?a��!���꜁cG��0ڇd)SZn��ᵢ� �|j^���BaW��NwV�j�N���/U�eW���o��_�ےRHƖ�`�����~�o`��X�Mqs~ע�;e�ޚ�-ʬ�M�ʐ� �� aU�2�$m-�ȇ�1�)���m�F�[��SV}�S����J�Y��0k|GD�^�R��r;��ϳ�������)�s��/�q�w*=9�y��(S/�E"��g�p���������J>'J~�����V��,�(�Z֍�8�?�:�5`�{S�xz~���OᏳ�o��p;��2ڜիe�6���F�w�^�ay�1��Ly�w���u�O���ѭ����3�(wM_c�i����sF��K�X�h��e���W�n�ً���B��z��5����G�1	/]K��h�HG�-�Km�->�,�����ӿ���U�ݗK� ��&�v�S�&�eM��=�zd=&yoJX�S~T���ӥڄ��qI���fۉM��Ҍ�b�!�y����늬�^ڛ�����q���c�~�����Z��W-`��xz�����{翡��z�̽�㍣�%��u��ӹ�O�~;�y��zz�@����<�������qzzJ��(n��;s���\H{��˨|�Ks�]�X�^C(�S���({��u�9=�{~���p�#p�Y�ݏ�fH��;;x��<^ނu>�}���qsvrr:��Vyj�;���8jv_�������gp<HϽf��m�Չe>�����X�Ҵ[��ӕK�)|��-��яE9��Ӛ;�~D����)����D��UF�c����=s�L�4KI���R�B:�����z�4K\@7G% #��������X���?��3��?��O����E�wI�N��{E�}�hɐK��x%2�1{�q�A'~����r`�i�([ߕ⋾cI�����.�C�p2���ow*��=��5It4W���g"	����Ɏ�'�������3�f�l`�5ڪ6B��GY�k���� ٔJq��lFQ�~�mn�'�w��+��˃�ª}j������ׅ��*k�	s!>�z^:)��C��0j�Vv�s�xL)�ˡ�|Q3yB_�o���z��5��Z���j+�5�O�w�=�-�3*F�P�X�_LlD�e��/o��/"W�s*V]l{S�v��,O%s>�◤B�؆Q{��ɉ*n��V���#� [ֻ���B,���~��*u�L7G�J*渭ݦ�V�*~�l����xp>ZJo͆����Kj�'8�N~���U]Q-xB.��Bm+�(�Jz�]n���>KP�2�ۉ���n?M�6�-��	��b�M�`kY���=���\}l�3�o^�O�+�ۢ�?M;@z���4ּ&[q�:~�kY^{�����ؽ������\:w/|���ԇ��7�f�A�үyڌ�3/�^�}p}bȴ����kq`�ʜ�k��&�.F�4�\IB��r��B�YIӮj�g�rMJ�́�-�Dǥ��#��_�N|���ɬ\<G�a��^xb�0�3wA��ޒ�+���oEk��>��O
�\����W��;�O@���n3rox7S��ݩ�\���g��~�ng�F����p ]�e�����8�ѱ.q�i��h�M��u�_X�r��$ަr�s�L���Sa���(s��;�ڈ����qn�%��з.f�]����mo�;�,_5�$��'�w����C'�������pl��mj� IB�R���tc��@��������H������t$τI_b-�̲c?�;�M�&�6!mF���rP�����}�2�H6(ұ	�����S-�U����	��@ELT��"�p�Ǒ\}�<�UׁY��i��c�24K��7�#�c!yL#�X?�D��8��R�+lJ��$M��A�XX4�?�%p�ruM�_,
����e5����j��1с�j�
����1|�Hd��>�9�%�a��/�]��P�I����reS�9 n��H�Ք�qAx��I�ҋ�X�<�$ɮ��3��o��`N���v=�u���L�m�0Ͽ�B6�۰�D�"7��@��W��x���ٰ>����c�Tx{��@ђ��x�.�ǛOvj]�L�V'�s1�UF[�i	�85�tyV�|��Gg�Ӟ�kO�%��^��	�����5Z�>S�3�,���H331��寐P�(�-�xF�y0�eAg�i���t���a��4��d.oǛ���� Ƈ⠚��X#��4���^�qĵ���1am�ʜ��U��J��Z'Q@7��s� �b��Ƶ�q�k��%��/��T�|�X�8�� GN�bE?5������ J+���ք�b_��:�ö<���a�<��cp ���OB�3��+��\6�S������5A�'Һ���o���zMXi��xWS�MpVK�b�4'qT���f�rJ-���@f��ʄ�OdJV�uQ�(m�WY�L4.X�<��_��rr慐[���U�lH1GZӠ2���aEj�u��!
��g$�L���4i0�~h�y=��Ҙ+f��J6�[v�����t��6�}B?Fl��'��I�H�Ns�+�h��}�-�24鵲p[=�l��e���҉�ӱK�z2�%QI�e��ԓ�yL4;��{3��^H��`E��TTJ��B�a+�i.�c6�ג��@,�QRF_-��jS��a+���\fJ"#%Š����MuF�OII��;�nI�CTc�(��Z�����-d{����ld�e�L�)l�����R��O̎���A�Q�g�Ыl�-X�v6�bb�� ��}T��UD���k�	���XW5�~�Pi�o��c!|�o��x��1�fg������&¥�a�f�n�����KDj��2��&�M� �[w
0U��
f�Q;�s$R�ϯ*	"�E��U%Ŕ��נ�(��0#fF`��!!o�+䊒�v�@x�?>�x��
@�_�u�1�ȿ kO��'[JM3�J��� �b���PK�:k[��҆��Z��$d�i��|:���p"-�%h'daeE�N�}C]L�DK�Tք�b��w��`�1���5�(���Hq�gG{1Z�F�.$q{��8��-WO-g3eެU�Z^��(#��`���p�����m)���k蟤6�ᩗD�H�e���G��tf�<���3���^��B�_�-�����w��r�[�b}ebCN��n�߾ϒTC����[��O�Y��l8Ri6Y���e�a��#*)���,�9�i����ǋ��x+����$��
�n�6P1��e��:I�-��\��N>ш^I���'�a�T�k��<�e��e����P�`�kO����!7"ل��9�����恞�c�t@�?�4��kK��uK��Υ�x�F��?Z�S�ʧB[meo�x����1nk�J����$j��K�v��{��}ň���&�<�X4c<����+�0�5�*�aV��o����v���t��5��娨�ZZ��\l�#\>�k��MQ�����ӧ���>�f�N �O������:m�$7�]�(��{�f���oawy�_/�o�v�)E�~r��YlJ���`ddljq$mz�����va�HYf�n�B@��r���t;8�����6��ї��&o��zBF��w�K.D��䤕��$L��PK   vm6Z�ւ&a  �     jsons/user_defined.json���n�0E%�SvU�dѪ�cUE`�Z%6��	����C�,��DbiϽ��#�����R������9�k#�����^ ;�+�Ԡ�m\<���;�����'��k�(󖯕���^���~�+	6ZƄ��r).��o�I�'a\�>)�=�&;Z�Vw�/K�M�EӎAOEy!�k�|��KY)���6�0M��w��ˢ �(�٩����b/"MF�ؚN��"�%{�� zh���^Զe{~�����`�s+���|�i�������&h�CWym.a�S��ؗ��	;�-7��g�M&l:;����zB���s���e�1�B�D��U�u+��R�+GpX?PK
   vm6Z&�@7  ��                   cirkitFile.jsonPK
   �V6Z��Y��k |l /             d  images/7c65d56f-74cd-491d-b8f1-3e526f205bd1.pngPK
   vm6Z�ւ&a  �               �| jsons/user_defined.jsonPK      �   ~   